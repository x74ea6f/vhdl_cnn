
library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.piping_pkg.all;

package fc1_rom is
    constant FC1_M: positive := 8*7*7;
    constant FC1_N: positive := 32;
    constant FC1_DTW: positive := 8;
    constant FC1_P: positive := 1;
    -- constant FC1_P: positive := 4;

    -- function intv_to_mem(intv: integer_vector; constant DTW: positive; constant P: positive) return mem_t;

    constant FC1_W_INT: integer_vector(0 to FC1_M*FC1_N-1) := (
-30,-6,-5,16,3,1,0,-23,-29,-17,-8,2,16,19,0,6,-2,-6,-12,11,7,-2,-1,13,6,3,-18,-28,8,12,-6,-19,-7,-22,-15,-12,1,-11,-16,21,-2,-4,-31,2,7,19,-1,5,-23,-2,4,-8,18,-13,19,-9,-6,-12,24,15,9,-11,-31,-25,5,-27,0,62,-11,-47,16,26,9,5,8,-16,8,7,0,12,4,-11,-4,25,16,2,-3,3,-17,6,-4,-24,0,5,32,12,-23,0,-36,1,12,3,-17,7,-1,-11,-4,2,6,21,3,15,-5,-17,-22,-34,12,23,4,5,30,16,-9,10,11,-17,-6,11,18,6,-17,-32,-34,-11,-12,-26,-7,-4,-2,-3,-20,1,8,5,16,5,-9,-9,-4,-24,9,-4,-13,-9,12,-33,-12,5,21,37,-10,6,-7,-38,1,46,83,-39,8,2,-11,-11,6,-19,-34,-5,5,-5,-8,-24,-12,-24,-17,5,-20,-7,5,18,-30,-3,19,7,-2,25,33,-29,-6,0,18,54,15,-38,-21,-17,-18,7,32,27,-67,-45,2,18,24,18,6,-97,-48,-11,-12,-8,-24,-35,8,29,4,-56,-45,-1,-13,2,33,6,3,7,6,21,27,6,3,2,33,14,15,19,6,-12,-23,-13,8,-16,8,-36,14,-3,16,23,30,7,-52,8,12,-13,10,56,24,-46,-3,15,37,-7,-24,-35,23,19,15,-11,-5,-25,-15,11,23,-1,10,-2,1,19,1,9,23,24,15,44,38,14,-30,7,12,6,25,17,8,10,-7,9,4,16,26,34,7,-19,-14,-14,13,5,-1,4,33,8,-12,26,-21,-34,32,24,28,-3,10,-35,-13,21,8,-3,-28,9,-1,22,12,4,9,16,-8,13,11,-30,-7,-3,-6,-2,-16,18,-7,-22,9,0,-19,-18,-7,11,-14,-1,-25,43,51,15,-6,20,-20,-42,30,38,55,17,31,16,-27,10,-10,7,11,20,2,-8,-54,-5,-9,20,20,-2,-1,6,-9,-24,
-27,26,5,18,-6,-11,20,10,0,12,-7,10,18,25,6,-10,22,-17,16,13,19,-15,4,-4,11,19,5,9,7,-5,-8,-23,-20,11,-8,7,15,1,13,18,14,14,-6,-10,-5,-9,-14,-18,-20,-26,21,25,22,6,7,-14,-6,7,41,18,-19,-35,-12,29,2,-18,18,16,18,-35,1,-1,-28,-23,11,-8,-17,-9,14,7,-4,-18,0,-49,1,-6,-9,7,2,-5,-15,10,-6,-9,-8,-20,0,-7,-19,-15,10,-11,-32,-15,13,6,11,3,17,6,1,42,-14,-16,-12,-20,8,-5,22,-22,-9,6,5,15,14,17,-12,6,-9,-9,4,0,6,-13,-3,-20,4,-4,2,2,-19,-13,-5,-15,-11,6,-4,-31,-2,21,-1,28,10,-29,19,11,5,43,24,14,-34,28,5,11,8,29,50,-38,-8,0,11,0,9,10,-30,6,26,12,-11,-3,19,-43,-15,-1,-5,-8,-1,13,-24,-14,19,4,4,4,10,-32,1,-41,-85,-73,-18,-29,10,12,-53,-65,-75,-70,-28,18,10,-54,-82,-78,-61,-49,-56,-8,-13,-27,-15,-14,-10,-50,0,13,4,38,-27,-52,-27,8,-22,-10,-14,-14,-25,3,25,-2,19,28,28,36,20,9,17,4,20,13,6,22,15,-10,22,28,-17,-61,-59,-4,-10,-11,-5,7,7,-51,-18,-21,-21,-2,-8,8,-48,-1,14,8,-5,16,14,-53,7,5,27,-11,-17,-12,5,9,20,4,21,29,8,18,7,21,7,-5,-18,8,22,-6,17,-9,2,29,19,6,-18,26,0,4,13,-13,-13,-15,31,-17,16,32,17,2,-21,12,-1,-16,-9,-9,-7,-3,-12,3,-6,-26,6,21,17,3,5,-11,-13,1,4,1,18,9,15,7,38,27,-10,14,16,32,22,25,10,-1,40,15,0,54,26,-78,4,29,0,-10,16,17,-40,14,2,-1,-24,8,15,-11,16,7,10,16,-14,2,6,12,18,-6,18,-3,4,12,
-4,-15,3,-12,-23,12,20,-11,-2,1,20,-11,-2,14,-2,9,0,16,5,22,14,17,-12,13,-23,6,5,1,14,-2,15,20,8,2,-16,-11,1,21,-2,20,20,-6,-14,10,-11,13,24,23,-23,5,-5,-6,1,-11,32,-9,-1,6,-10,9,-2,-24,-65,-8,17,18,27,9,1,-23,-17,13,30,23,7,-23,4,6,18,25,-10,12,15,75,8,1,8,-4,-14,-2,-2,9,-15,-17,3,-1,15,7,-8,26,2,-6,-20,-13,2,3,-2,3,0,-19,13,24,-4,-7,19,29,22,25,-3,20,31,3,-20,12,-2,4,2,7,2,0,-11,-8,-5,-14,1,-1,-2,-10,38,3,30,10,-10,3,27,-8,3,-12,-11,19,-6,3,-13,-8,-9,-20,-6,-14,25,38,-5,-4,7,-13,26,11,58,-11,4,1,-31,19,-3,2,-24,-10,10,-3,-8,-8,-28,24,0,9,15,6,-4,18,-3,6,2,-13,1,9,-2,14,-9,31,63,50,45,-8,7,8,33,48,20,-12,-62,-32,-14,41,37,44,-13,-41,-53,-8,-27,-28,-12,-35,-44,-3,2,-24,-34,-42,-32,7,36,3,11,-2,20,10,45,34,30,29,1,3,34,1,-18,-7,-12,19,-28,-17,22,-45,-3,-10,15,16,-4,-10,-99,-7,2,-5,24,-33,-28,-41,7,25,-22,0,-28,-21,-27,-5,-30,-40,-37,-27,-13,47,15,-9,-8,-12,-25,18,39,14,6,9,-8,15,23,-2,-13,-6,-6,7,-5,13,-3,-9,-23,-5,-4,-19,3,6,0,-16,1,14,0,-1,-19,-3,-3,0,3,8,1,-23,19,14,21,6,-8,21,-13,1,-3,17,-8,2,4,17,30,31,-13,-21,12,-11,-18,-6,-13,23,-7,-12,20,-45,-6,-41,-21,-18,-27,-6,-69,-15,5,-8,28,35,35,36,-8,13,7,22,6,64,69,-14,26,31,45,-2,-5,48,0,20,27,-4,-31,-10,50,33,34,17,6,-33,-33,40,
11,-6,-21,-15,18,-5,12,11,0,11,-10,-13,-20,-4,-15,-3,16,-18,-23,17,2,-6,-25,-12,18,5,11,0,-4,0,20,7,19,2,-19,-8,-8,26,-1,-8,1,3,-7,13,13,27,26,44,29,1,12,-1,-19,-2,20,25,-14,22,24,-13,-13,4,24,17,18,18,-4,11,2,23,33,8,12,-9,16,-28,-2,27,0,-25,22,-2,-10,43,-16,11,-3,1,42,20,17,-7,-7,10,13,14,14,42,35,20,22,11,10,30,23,-4,-11,-10,24,-2,0,-15,-15,4,-16,7,17,15,27,9,-19,15,27,-7,-2,11,9,-11,30,-1,10,-5,0,-9,21,49,3,18,2,10,-10,-9,8,3,-3,9,37,19,28,-19,2,-6,-1,31,9,4,0,-40,-60,-50,9,13,-18,9,-7,-35,-16,58,15,17,6,-28,12,29,61,-4,-10,14,3,14,-7,40,13,17,-13,-23,-26,-1,11,8,-7,-1,-18,-30,1,18,27,67,27,56,-5,46,27,-13,-54,-14,61,125,80,0,-24,-18,15,59,93,70,33,4,-12,-17,13,38,-7,6,-5,9,2,5,15,-4,7,11,7,47,42,46,5,-10,-27,0,29,13,7,2,13,9,22,-4,5,22,-12,4,-14,8,2,-14,-18,-17,42,-4,-22,-6,35,34,21,48,3,13,-1,2,18,-12,26,17,7,-1,27,25,-3,38,11,20,12,12,37,3,-16,-19,-17,38,-7,-8,-5,18,-14,3,-3,14,27,15,14,-3,-5,-10,22,0,6,-1,-13,23,-7,-2,-12,3,28,9,21,5,17,5,-1,18,2,3,7,-12,25,-5,7,-3,-2,12,21,10,13,29,-25,-34,19,31,20,44,33,0,2,6,-12,14,-19,0,-8,24,-10,-4,-78,-49,-15,0,6,0,-43,-67,-42,26,25,11,8,-46,8,6,33,11,5,-18,-30,14,4,23,12,-4,-27,-16,-26,31,13,-7,-11,2,-52,-51,6,-5,
8,13,14,21,-3,-35,2,-4,5,19,-5,-5,18,15,3,8,-1,7,-6,-9,-9,5,18,5,4,30,22,9,-18,1,-9,-25,6,8,5,14,-5,-1,15,-12,-13,12,17,8,-12,-26,-32,-6,9,-25,14,25,2,3,-2,-23,5,8,33,-5,23,24,60,9,3,-56,-28,5,29,3,24,-1,-30,3,8,2,-30,-8,10,-1,28,-37,3,-47,2,18,18,-1,-6,13,5,-1,10,5,5,6,-8,0,-21,-28,-29,-29,-4,-24,-5,4,5,-7,9,11,15,7,-18,12,16,-14,15,24,15,-14,22,11,5,12,17,6,-5,21,4,-18,6,2,1,-11,-19,-24,-11,-13,-11,2,4,-11,-11,-2,-21,4,4,-12,24,-1,-6,34,17,14,-4,28,36,-10,-36,-46,6,29,7,31,9,14,-4,-23,-10,7,28,16,30,11,7,-9,30,14,29,-1,-7,-28,-15,2,5,6,-6,18,-13,24,3,24,16,-2,20,-11,-7,-93,-89,-55,-52,-30,-20,-27,-30,-34,13,23,86,47,-21,-38,-39,-33,15,1,0,23,-15,-8,-8,0,-22,1,7,13,34,29,18,-4,-45,-19,-31,-6,-32,-46,-41,-5,3,-22,-1,7,-7,-12,30,-28,1,4,20,36,-2,46,-24,-8,28,-17,11,-8,83,22,4,-39,-7,24,38,-13,16,7,28,18,6,8,-12,-8,21,30,-10,-13,0,-64,-12,-19,27,4,-6,10,-28,-17,-23,-33,-4,-18,8,9,-36,-14,-4,-16,-8,-36,8,-42,3,26,6,3,4,27,3,35,34,-19,18,19,31,5,5,-10,8,13,18,-12,-11,15,17,6,21,-8,-7,-29,-4,-25,-10,-37,-12,8,5,1,21,15,-10,1,-6,-55,-1,-5,-3,2,-20,27,-7,20,21,5,-9,-1,61,-5,30,27,-15,2,-6,-25,6,18,-41,-16,11,-1,-78,-14,28,11,-2,30,9,-31,-1,4,19,1,33,-5,-30,-10,7,23,64,56,8,-20,
-6,-15,-16,27,-15,21,3,-19,-20,-4,25,26,10,14,19,19,-12,25,14,-5,-8,12,9,-17,29,26,-18,-7,1,9,-18,-8,12,21,6,8,32,5,-3,-4,3,28,2,18,-3,7,3,-6,-1,7,-11,-9,0,-10,2,-5,14,11,6,30,4,-33,-14,11,-12,9,50,43,11,-35,-21,-28,-8,-13,-34,3,28,-1,-15,27,-22,-8,2,-53,3,21,1,0,-4,14,13,5,11,44,38,31,-5,-14,8,4,0,24,-8,-1,-4,-21,-6,18,32,24,8,-7,33,12,4,19,24,26,1,7,-14,-32,18,-3,1,-2,17,-15,-13,8,7,1,7,7,9,4,-6,4,25,15,4,5,-1,18,15,8,-16,11,-19,7,-13,-9,-31,-15,-19,-10,-14,-13,-17,-41,5,0,-11,-10,21,2,21,-30,-14,-11,-6,9,-21,-23,-23,-4,-5,1,-13,8,-4,-38,28,-5,-10,-9,26,10,5,-2,-2,16,5,1,-3,-7,13,-38,18,11,-13,-53,-18,11,-4,89,29,-57,-67,-38,13,25,105,64,-43,-56,-35,6,26,49,23,1,22,1,17,-26,-5,8,-38,-53,-42,10,15,-12,-20,-3,18,40,3,20,10,-14,-21,-20,-3,5,-36,-6,-29,-13,-14,-35,29,1,19,41,15,-35,-40,-2,-22,13,93,27,12,-31,8,-4,15,12,-41,-12,39,-5,-18,11,15,-20,-40,-52,37,4,13,1,10,7,9,11,6,13,34,10,-2,-3,26,-19,2,-14,0,-5,-10,-10,-16,-11,11,16,-5,-17,19,10,-19,44,27,15,-3,15,-36,-25,36,-23,-14,-14,-1,-5,-17,8,-42,-10,14,11,30,-12,-23,3,8,15,18,10,8,26,10,7,-28,15,-14,1,-1,-27,-24,-12,-7,-20,-14,-20,-28,-58,-6,22,-6,-46,-7,22,-9,27,2,-40,-2,15,-29,-3,17,-17,-3,-14,-22,-27,-16,-15,26,-9,20,19,-23,27,4,24,1,15,17,17,16,-15,
0,11,-8,11,4,26,26,-21,-2,6,9,-23,-3,19,-4,13,-17,-32,-20,-11,-4,-2,6,5,54,2,-13,-18,-18,6,15,10,1,-4,-11,-25,-7,-4,-3,1,-20,-12,-17,-9,-15,7,-5,7,-9,-12,40,13,16,22,25,8,-14,13,21,14,-22,7,-4,16,-8,-17,-21,26,19,-29,0,3,18,-11,1,-4,-14,1,19,-11,9,20,-12,-5,-3,10,-12,13,9,10,-28,-30,-24,0,-9,-11,4,6,-1,36,44,29,17,29,22,-22,-7,-11,9,16,-10,-8,-5,8,-28,-13,-26,3,24,5,-15,2,35,23,25,2,5,21,39,3,19,-15,3,0,-9,21,10,26,-24,-1,-28,-30,-3,18,-2,14,10,-21,43,6,13,32,7,7,-6,1,-1,-7,-19,-56,-1,3,18,-18,-22,9,-1,-17,7,13,35,-9,-45,-3,-17,15,25,31,15,20,9,-10,6,-5,22,-7,-12,-9,-22,-10,-22,17,10,-1,4,-15,37,30,-20,-34,10,-2,36,-26,-60,-92,-10,47,65,41,17,-33,-39,-78,11,36,-9,10,9,-38,-57,15,17,3,-18,-1,1,72,11,7,-20,-13,-26,18,29,17,-25,4,-29,-23,4,-3,14,0,36,-17,19,-4,31,38,-1,27,-17,39,36,12,-32,-23,-10,22,-27,-20,4,22,60,8,-19,26,14,13,-28,17,-29,-17,-2,33,31,48,-5,-20,-44,-2,50,27,23,-5,-25,-33,-13,4,0,-8,-2,17,-23,43,41,14,40,13,32,-21,12,-6,1,-4,10,8,-19,25,-6,-44,-14,14,9,-20,15,0,51,43,26,-4,-20,16,27,10,2,-24,-12,-39,-10,-5,0,29,-11,-7,-30,-30,-14,-5,-15,16,-14,-9,31,7,7,52,7,1,-32,15,9,5,-41,-35,-3,-1,14,27,-7,-23,-51,-52,-15,0,-1,-11,-29,-28,-54,-20,13,15,-30,-10,4,-16,-14,14,-15,-12,-4,12,-52,-36,-18,-31,-43,-25,-4,-18,
13,-12,-13,30,16,-10,16,8,5,10,-26,-4,1,-21,16,6,-1,-12,-22,-18,4,-10,11,2,42,1,-11,12,12,-3,-6,26,17,7,-6,-5,20,14,-1,30,22,-5,-18,-39,-16,-1,-6,-21,-14,15,2,17,29,17,8,13,12,-2,6,-11,5,18,-3,-6,-16,-11,-12,-14,5,48,1,-2,33,6,-9,37,41,-6,5,31,-8,13,15,24,12,2,-3,15,0,-4,-4,-31,-32,-35,-16,13,10,10,1,1,15,33,30,31,14,11,5,-13,-9,-23,-11,10,-1,-21,-34,-32,-28,-8,-24,15,29,0,11,10,-16,-14,-3,20,8,30,-5,12,11,-3,-14,-27,12,22,31,0,-32,-11,-15,-15,-22,0,4,-3,-8,18,39,27,46,-6,20,12,27,49,26,38,1,15,7,7,-11,29,-15,-5,-11,-11,18,-6,-24,-42,-19,21,-12,23,23,-13,-4,20,-7,-2,-10,0,25,21,0,-2,-14,0,14,2,5,-19,-8,-16,-9,-8,9,-22,-23,-11,31,6,-71,-37,28,55,14,21,-21,-76,-88,-9,31,11,-1,28,-18,-2,71,49,19,-2,-24,32,29,48,45,-8,4,-21,6,35,65,34,-25,-5,10,-2,38,38,-22,-7,-4,9,9,13,12,47,-9,-8,-14,-16,12,25,34,-16,-20,1,-42,-20,-28,61,-12,30,52,-1,-39,21,43,-7,8,12,15,20,35,90,-3,4,3,0,22,45,40,-39,-12,-19,-7,20,36,-12,-13,29,32,23,31,38,21,16,-12,-6,0,-1,-16,11,-1,-12,-3,-28,-13,-3,5,-4,1,17,30,-24,4,15,-4,24,23,5,-7,24,10,-2,-10,-23,-29,-2,10,10,-38,-33,-39,-15,-32,-33,-35,10,39,19,65,36,31,68,10,14,40,42,65,63,54,-19,-10,-17,0,57,33,21,-1,18,7,44,-14,-30,34,-5,15,58,16,-52,-32,-16,1,-2,16,7,-13,0,-7,-29,-32,-39,-11,-20,-24,23,
-4,8,7,-4,-16,-12,14,-7,-3,9,-9,-1,-19,19,-13,-6,25,1,19,4,-18,-18,-19,17,3,31,24,-19,-1,3,-2,28,16,-12,-17,-16,-13,4,-25,-23,-10,10,-4,41,16,-18,0,5,-6,4,20,14,-8,-4,20,20,22,-14,-4,4,4,-3,-3,0,12,-8,20,20,-10,8,-9,1,-21,32,6,-40,15,-14,-3,2,36,-39,2,-8,-5,-2,12,4,-58,3,7,12,22,17,36,-6,-4,-2,-5,-28,-43,-28,-39,-41,-9,25,3,-4,-10,1,-4,33,-28,-33,-3,16,-1,-12,-18,-18,-10,6,12,39,13,-21,-25,12,0,17,9,2,-12,-11,-19,-7,3,-33,-32,-5,25,14,13,-6,-14,13,13,5,16,-15,-26,0,17,11,-5,-20,26,48,38,42,1,-2,12,12,11,5,40,-7,-28,5,0,12,12,-3,-7,-15,13,23,37,-32,-3,-8,2,-3,8,-11,9,-5,-12,11,19,7,18,24,12,-10,-19,-62,-26,-35,-12,-56,-28,17,45,17,-27,-87,-73,-6,2,-59,-92,-63,-74,-63,-36,-21,-18,-26,22,-61,-58,-30,-16,22,49,20,41,3,-7,-34,-21,-42,-10,-30,-51,0,2,14,-24,-43,-21,16,20,2,5,-9,-5,-30,-5,10,2,-20,15,2,4,-39,-29,-6,-2,-5,-10,-26,-36,-36,1,-2,-3,14,0,-36,-13,-22,-7,-1,11,-44,13,-6,-16,11,-30,-37,-21,-11,-6,22,-18,-11,-28,-20,16,12,4,6,-8,-14,-25,-30,-9,7,1,2,-1,8,-9,2,-8,-11,15,3,34,-37,-24,-26,6,2,14,28,-11,-16,-17,-5,-15,13,-1,-30,-21,1,-21,-18,1,-34,-8,-13,14,38,8,-32,4,-1,18,-1,1,-12,-12,-18,38,-16,-2,-10,11,38,38,39,-24,-7,-8,8,57,63,44,-43,-21,22,9,18,38,7,-17,11,8,-8,27,-6,-16,15,1,-17,26,42,0,-33,24,26,40,46,71,58,14,36,
7,-21,-31,-17,-3,32,20,-5,-2,-16,11,-8,15,12,6,3,-6,-12,31,14,26,24,-21,8,-1,3,13,11,-13,-4,4,20,-12,-21,-18,-22,-19,-5,-20,-4,6,-4,-19,2,9,6,31,33,-14,2,-16,-21,-34,-17,27,-4,8,0,5,16,-12,-11,-59,-13,11,24,37,30,3,-16,10,-7,1,29,21,-27,6,0,-3,-9,12,23,-16,38,-2,-16,-14,0,13,4,1,14,30,29,18,-11,-9,-1,-1,33,36,4,27,28,21,-11,-29,-15,23,2,-3,29,-2,-3,-3,7,5,11,3,18,-26,-16,33,14,29,-18,32,9,-4,0,6,2,13,16,5,6,0,20,-1,-4,-1,5,21,1,9,0,3,25,1,-12,-34,-20,-50,-4,-11,-1,-43,-45,-13,2,-12,-1,-27,-14,19,-6,6,10,17,-10,-35,-11,-14,0,18,-4,-11,-6,-13,-16,0,8,-20,-7,-6,-17,-19,-19,13,-2,16,-13,-20,-20,-24,7,2,69,74,61,22,40,21,3,17,29,45,36,-67,-64,8,35,44,34,17,-4,-35,-17,12,7,18,19,-20,2,0,7,31,16,-4,1,11,17,-8,27,26,22,6,1,-6,10,-17,-38,-23,-4,12,30,-20,-27,2,-24,-2,-59,20,17,33,24,3,-1,-123,-2,15,34,52,16,-5,-27,-6,-8,-6,14,-5,-8,24,-5,-12,6,20,27,-8,14,22,31,15,4,8,0,-4,-17,0,-3,-10,-31,-7,13,11,1,13,-3,-2,18,19,18,0,-6,13,3,-19,-30,-5,-20,-12,22,-8,-18,-17,-10,-13,-10,29,23,-13,4,8,-15,-12,17,20,-12,-1,29,-17,9,2,-1,6,7,-4,3,22,-1,20,30,28,19,11,-22,-15,-20,-22,-56,4,5,-19,-39,-63,-57,-115,2,-11,-19,16,-7,-36,12,0,-13,8,-12,-7,-4,68,12,-30,-44,-24,-5,5,13,16,-4,-13,-26,-16,-10,-13,-22,-7,15,-15,1,-13,10,
-9,11,3,-1,-13,-12,-13,3,-6,9,12,9,1,-9,-7,-7,-8,-7,-16,8,10,-7,-5,4,-17,-6,-20,-16,-8,13,-13,-5,-20,-3,-3,-3,12,-8,-18,-14,-7,-4,-15,-13,14,-10,-19,-7,8,14,9,-15,12,-17,5,-6,-18,-19,-2,6,-7,-5,-8,13,-11,7,-14,1,-3,10,-3,1,3,-19,-17,-2,12,5,9,-13,-14,10,1,-19,2,-18,-12,-15,-5,11,9,-9,-20,-8,12,-16,-12,-7,-15,-17,-15,11,-5,-10,9,-19,-16,-1,-15,-4,-2,-2,12,-13,12,9,-17,1,-16,-20,-7,11,-11,-1,8,-19,-5,-13,-19,13,14,14,7,13,13,12,5,-18,10,15,-3,-5,-18,-18,-9,6,-5,-3,-17,5,8,9,0,6,-7,-19,-9,3,-6,-19,-5,5,-4,-6,9,15,0,-17,-7,-1,0,-18,-14,-16,3,6,-16,11,-7,-6,-17,7,11,-19,-19,7,-19,10,-15,14,-15,7,-3,-10,8,-18,3,17,-11,17,1,14,4,2,-16,-17,5,16,1,2,-14,-3,7,3,6,-2,-1,-7,-7,-7,2,-3,13,13,2,11,-2,-12,4,-5,15,6,3,-5,5,-7,-12,-2,-13,-1,11,8,-8,5,-1,-6,16,8,6,-8,-7,-14,-7,-1,7,10,8,13,-8,-17,16,1,-2,14,6,7,-13,-14,10,-2,-5,-14,-6,-3,9,-11,12,-4,0,-5,11,5,6,-15,6,2,-5,-9,-8,14,-7,-18,11,-9,-7,-6,-3,-11,-17,-19,-8,-11,-4,-7,4,6,-14,-5,0,-15,-10,-15,10,0,16,10,3,-19,-10,-4,4,-16,-7,5,4,-1,10,-14,-3,11,9,-18,9,-15,-16,15,-7,-13,5,12,-1,4,-7,13,10,-17,3,-17,16,8,2,7,1,12,-13,-2,11,-10,-1,-10,-16,-19,14,-17,10,-6,-7,10,-5,-17,14,0,0,1,13,-10,8,-1,-10,5,3,-14,-4,-2,-16,-1,8,12,-13,-8,-1,-5,
8,5,2,-8,11,11,17,19,29,28,9,15,14,0,0,28,-10,-14,-10,13,0,-12,-7,-10,9,-4,14,14,5,18,-8,26,3,11,-10,16,10,-1,23,24,-7,-37,-3,-8,10,23,21,4,-8,10,-16,-1,3,9,13,-6,15,4,-5,-10,-1,-16,-39,-29,-26,12,39,6,-22,55,3,9,73,7,-25,12,33,9,-5,26,-8,24,-11,74,16,-6,6,-12,-18,1,1,-14,-40,-20,-24,-23,-15,-12,-5,36,5,36,15,3,3,8,7,17,7,-9,20,9,0,11,-12,5,-5,5,-14,-15,8,-29,-2,-15,-7,-11,-6,-10,28,34,2,21,-6,18,-2,-14,11,-2,9,-36,6,-23,2,-13,11,-24,-36,27,2,15,1,-12,5,-12,20,22,-13,12,39,26,12,-21,-25,-39,20,14,-19,12,-21,-33,10,10,-15,-36,2,-6,6,23,-5,-43,-26,38,19,-14,19,8,-5,7,12,16,-16,-9,7,9,-18,-9,-14,66,62,45,35,22,7,5,104,62,-17,-27,-90,-25,16,101,94,36,-23,-19,0,-39,-5,-37,-66,-40,43,37,-6,-30,6,3,40,90,59,26,9,11,7,39,64,-1,10,-3,-6,2,24,1,-49,29,-8,4,-4,-1,7,-23,-6,5,-42,-3,21,5,-59,-34,-2,11,-4,-39,-46,3,-5,6,27,4,-38,-7,54,-13,-39,-12,-22,-14,9,91,30,22,8,-3,-4,7,4,-2,-10,0,-19,6,11,-41,20,1,-2,6,20,10,4,6,-6,13,16,-15,-9,-52,-32,-25,-31,5,-9,-22,-30,-41,-15,-7,42,-38,-30,1,12,17,20,28,-5,23,9,11,15,1,-3,12,0,-25,-10,-2,-26,-9,-18,-42,-8,16,-6,11,11,5,35,-22,1,-8,3,16,42,25,-18,-27,-9,-67,10,46,8,66,-32,-43,13,36,-11,-32,66,-3,-3,43,7,-82,-25,5,22,5,21,-7,-51,-40,48,-11,-6,-12,-32,-49,-28,15,
-20,-4,8,11,30,0,-3,-15,18,5,28,32,15,10,-19,4,2,20,14,-18,6,-4,-6,-1,25,-2,6,8,-14,25,-15,10,13,-2,8,-8,20,-1,8,16,7,12,-6,5,25,27,-3,-20,19,-2,-11,-17,5,-3,5,12,-7,5,23,29,21,7,38,12,-3,-16,-9,25,14,32,-7,-39,0,2,-8,-1,61,27,-2,-3,9,-23,17,-35,24,9,19,16,21,11,11,7,12,27,24,21,-17,7,12,-11,-11,28,29,-13,-18,-37,14,26,39,32,11,10,-12,8,-25,-14,-2,-9,19,-1,-4,5,22,5,-2,-16,3,4,6,26,15,-2,-11,22,12,15,-15,13,-3,31,-2,3,25,14,-7,5,27,-24,-1,-1,35,16,-19,17,-24,7,13,17,-19,-23,12,-1,-16,0,12,8,-16,-3,-8,-8,48,-15,-42,-26,8,-1,7,10,3,-2,19,-7,11,-1,-9,25,13,19,18,-27,14,7,-10,-1,-3,-5,-33,-54,0,-40,-42,-12,-27,-22,-19,35,16,-5,-5,-4,5,-26,21,-26,-7,9,32,-20,42,69,38,41,24,41,5,0,33,68,3,-31,-66,10,30,0,-34,-3,1,-7,-10,3,15,27,14,-5,14,-15,-8,22,30,24,8,54,-22,4,25,41,32,2,98,0,-15,7,43,35,20,55,-11,6,28,31,-40,-18,70,6,7,52,53,15,11,-60,-12,-18,11,42,16,29,3,0,20,31,14,23,1,22,-24,-35,3,7,-5,19,18,-14,4,11,23,42,27,24,-9,15,-9,-4,4,-14,9,-25,-34,-6,20,6,-12,-13,-23,-6,20,-13,-1,-13,-6,19,29,12,11,10,23,19,4,10,2,21,-8,29,-8,-1,-8,-16,18,23,-7,37,-9,1,9,2,25,-11,81,-10,2,-24,-27,5,7,44,-27,-32,-7,-10,-22,-45,-15,16,-24,3,-42,-20,-35,-41,15,27,-22,7,40,22,-27,-8,-1,22,7,23,33,-8,
4,-16,-6,-15,8,-6,-18,14,1,-16,0,-5,-17,2,5,-6,-12,-7,-10,7,-5,-12,0,-13,-16,-10,-5,-14,3,-14,9,7,-15,6,7,0,6,-15,-5,-6,-1,-8,11,-8,16,14,-12,-2,7,10,-4,9,0,-16,-9,0,9,16,-2,-17,1,-16,16,6,13,4,-4,-1,-17,12,12,-9,3,-18,1,5,7,12,-9,-9,2,-14,3,1,1,9,-14,3,-11,7,-14,5,-7,-12,10,-12,14,13,-1,17,5,11,0,12,5,1,-1,15,14,-17,12,11,10,0,4,4,-7,15,-18,4,-7,-4,-3,11,-14,14,-5,-1,6,-12,-12,-18,-2,1,13,9,14,-11,-16,0,1,-1,2,5,6,-13,-4,-6,6,-14,14,-5,-6,-6,-16,8,-8,5,17,-2,-16,8,-8,4,-13,15,4,-9,0,-8,-7,14,-14,14,-2,6,1,-10,4,6,-3,-3,-1,16,-13,1,17,-2,-18,-14,9,-1,5,6,3,-15,1,10,4,-16,16,-2,2,-14,-6,12,-13,13,14,-13,-2,17,-8,-5,-13,5,-7,-6,14,10,8,-4,-8,-2,1,2,-13,-1,-15,-15,9,1,16,-13,11,-16,-8,6,-1,7,-9,8,-4,-8,-9,-4,-16,-4,0,-8,14,-17,2,-7,-17,8,1,14,-15,9,-3,-6,15,-3,-13,12,9,14,-14,7,-14,-7,11,-10,2,1,-10,-18,0,14,-17,10,-14,-11,-17,7,7,-2,16,5,3,0,12,6,12,-15,1,-1,-15,-1,12,13,12,-16,-10,5,-17,-11,-17,-11,1,8,9,-7,5,-5,6,-12,-12,-16,11,-5,-14,-9,-4,8,3,8,14,11,-2,-17,1,-5,17,14,-2,6,0,15,-4,9,-11,2,-13,3,-11,-1,14,-6,7,15,-2,9,-5,11,-4,-9,2,3,-11,3,2,-13,-13,-10,-15,-6,4,-5,-9,4,-1,8,12,-4,-14,-6,-14,-11,4,0,9,6,-6,16,-16,-17,10,-14,-1,4,
15,11,5,10,0,-14,-6,3,-12,-2,-13,4,-5,-24,19,-2,-7,0,-9,2,-10,-5,15,26,-10,-5,17,8,-11,10,18,-1,12,2,10,16,-8,-14,9,-17,-18,11,3,1,-6,-9,-21,-18,24,11,10,10,-14,-3,9,-11,-25,3,5,-12,1,-12,-25,-5,9,11,-27,-5,-43,-12,23,40,23,8,9,-18,21,13,17,-5,19,5,-4,57,7,7,-19,18,11,2,19,-28,-15,-28,-9,-18,-5,30,-5,19,33,-11,4,-4,-8,-2,-13,-22,5,11,-1,0,8,-12,6,-26,-8,2,-5,12,15,2,-35,-7,-4,-8,-11,17,27,1,12,-11,14,-3,-2,18,15,15,6,7,0,-33,-2,-22,-23,3,25,18,10,-11,5,24,30,-3,-7,-28,-4,21,1,26,17,-17,-23,7,19,33,-4,17,18,-1,-4,-12,39,-5,9,22,5,0,9,-8,5,51,-8,7,11,14,30,34,1,13,-12,-15,-17,0,11,10,-32,8,32,47,8,14,-22,-5,27,12,13,2,16,1,-23,-16,-44,4,23,-48,-13,-16,-36,-50,-71,-60,-46,-12,5,28,22,45,29,26,32,-20,-5,18,14,26,40,26,-6,-11,-2,0,-17,16,24,11,24,1,-9,-6,-35,7,-17,-10,-18,9,8,-17,20,-6,6,-3,-44,-19,-3,1,-2,20,19,-6,9,-9,11,13,-12,13,1,-8,1,73,4,10,1,18,20,1,0,16,-28,6,-36,17,16,37,-1,5,8,13,3,-31,7,-11,-13,-9,16,8,-13,-13,-33,4,-3,-37,-15,-22,-1,10,17,26,-7,11,-8,-4,29,10,13,26,12,15,11,3,-9,-8,-16,7,-7,10,-1,-22,-15,-29,-41,-8,22,-3,24,-6,-10,1,-6,25,-6,-30,5,10,22,24,11,-9,9,31,6,1,21,28,16,35,34,-12,53,-4,77,34,6,2,-3,19,1,20,-20,-9,-22,4,-14,4,-4,0,-15,-47,-30,-8,-18,4,
-5,-7,-12,-12,-10,-11,3,-21,13,-12,7,16,17,4,14,-6,0,36,18,36,-10,12,-3,16,-35,-11,-13,-6,-3,-8,2,-6,-18,-8,-14,9,-1,-8,-2,-15,0,19,28,6,-11,47,60,-8,-21,-14,10,-18,-6,-8,14,-5,-12,-27,-12,-6,12,18,-27,4,-1,39,11,-20,-19,-22,6,25,18,-28,8,-30,-68,11,1,6,-19,14,-14,-67,24,-20,4,19,6,4,-6,-2,-15,25,15,16,-6,-3,8,-13,-16,-17,-20,15,25,-9,-1,-32,-15,26,0,7,16,9,2,55,39,13,18,-4,3,15,-14,-25,-14,-13,-24,-15,2,-18,-44,-26,-28,9,-10,15,20,-11,-11,7,29,5,26,23,15,-6,-21,3,-13,-13,-25,23,5,-3,-19,9,-12,-17,-6,-13,-2,-20,11,-1,28,8,4,13,-6,0,0,7,31,26,17,-14,28,-13,1,30,20,9,10,11,20,-11,-40,-5,-12,22,-11,5,22,-19,-38,1,-2,11,-40,-23,-11,-2,21,7,-55,-67,-56,-11,12,-8,-23,-23,-42,40,91,88,-19,-7,-8,-76,-20,21,-1,-44,3,-25,-57,-76,-70,-80,-51,-3,-1,8,7,0,-29,-23,34,8,31,37,6,-14,-22,-17,-9,1,-1,6,-8,-42,1,-3,-27,12,-33,-10,-33,-15,-7,13,7,-29,-19,-29,7,21,-5,-35,33,-7,-61,-19,-11,-47,-38,-16,-19,-71,27,3,15,-1,-28,-40,-16,15,18,21,51,-14,-21,-16,4,6,-22,3,1,10,-22,-2,-27,-7,22,17,18,-16,9,2,-3,18,6,25,5,-16,-6,21,-19,-23,-7,-11,4,-3,0,-17,-20,-22,-2,14,14,22,18,21,-15,-2,26,-18,-4,19,13,-33,-38,-2,-18,0,-14,10,12,-34,-31,-16,-28,17,-6,-26,-32,-26,7,-6,33,-24,-25,-39,-2,30,29,19,-1,-9,-16,7,16,35,0,17,40,-6,26,17,2,13,34,16,28,20,-13,11,-11,-44,-41,5,
11,26,18,-6,18,6,0,17,33,-8,-12,2,-7,-12,3,-2,15,-17,-11,-11,-3,10,-8,11,-32,-10,35,3,14,-13,-4,-11,9,22,27,3,-7,19,14,2,-9,22,37,19,1,3,-20,-21,19,0,30,24,5,0,14,26,-1,-14,-19,-21,34,17,13,-8,19,1,-13,-30,-2,14,4,35,-10,-13,28,3,-35,-5,22,-12,25,3,18,-40,-7,6,-4,3,11,-9,2,-3,-18,-9,-49,-20,10,39,-7,10,8,-8,-2,13,3,39,42,20,-19,-6,9,8,-26,6,38,7,12,1,3,7,24,24,-30,-20,26,23,29,-13,-8,-37,25,4,20,-8,16,35,19,-7,-10,16,12,2,-7,-17,-19,7,9,14,27,7,27,12,28,17,6,37,33,0,0,18,17,-8,17,44,9,-9,-18,13,31,30,11,11,44,22,1,30,3,26,4,30,30,-9,23,7,5,-2,-5,-26,20,26,3,18,-3,-1,-14,20,1,16,-45,-32,9,4,26,11,-21,-50,-30,4,57,31,-9,-41,-106,-7,16,46,39,1,-10,-59,-40,31,-11,-38,12,19,-20,-63,14,17,-15,-28,-13,38,32,0,-44,-42,-10,-24,8,1,-14,-11,-19,19,8,15,36,23,-3,30,-27,12,-28,-28,-22,19,29,11,19,-11,-47,-16,-1,24,5,-11,-28,-32,58,14,-56,16,11,3,-17,26,31,-23,2,5,20,15,-2,-27,-41,-15,-10,13,-2,-24,-14,-5,-5,20,-4,14,13,-19,30,-13,24,-2,2,17,6,-3,4,9,18,-16,-3,20,26,11,10,10,-55,2,15,3,23,-7,9,-9,40,12,-4,-20,-27,13,34,-2,-16,-22,-10,-2,-17,-15,-5,-7,24,-18,20,30,40,34,-4,0,15,39,26,35,27,34,-12,-5,-6,28,0,-4,-6,-79,16,28,29,12,37,1,-64,28,14,1,39,13,29,13,3,-9,-15,-16,22,-3,19,11,-15,-19,-30,-43,-20,1,
28,7,5,23,0,-1,-10,19,9,2,12,-4,-9,-9,12,17,11,13,-9,4,18,29,0,6,10,24,5,14,29,36,-12,12,19,11,16,5,-8,12,-8,17,23,8,28,6,21,14,15,43,39,32,1,2,4,24,11,27,10,-8,7,3,5,28,40,-7,-20,8,-21,-19,-16,84,20,-26,2,13,-4,-11,18,14,-4,24,12,3,-10,51,-11,-10,3,1,-7,20,14,2,36,35,46,26,15,6,42,-30,-13,-1,1,-7,6,31,-8,1,-15,4,-18,1,-18,-3,20,9,6,-7,6,-5,-4,-15,10,30,-11,10,33,-7,-4,25,12,13,6,21,23,21,14,-6,26,20,39,24,11,0,19,23,28,35,12,24,3,-13,8,31,24,28,31,-8,-12,14,30,-4,10,33,-13,-28,-56,36,7,-13,-4,27,42,17,63,0,-14,-11,22,-2,-2,24,-4,-14,18,38,44,30,47,32,18,-9,30,50,39,37,0,-41,-23,-25,-20,-4,-23,16,-5,-22,11,14,15,-2,-35,-10,14,56,22,36,66,9,45,32,40,31,-9,31,22,40,56,12,1,-17,-28,6,29,-11,3,-33,-6,0,5,3,-37,-33,0,-18,4,-26,-1,-16,-30,9,-4,-5,-10,-5,-17,-22,15,5,50,-16,14,-6,-14,-46,-2,41,-11,-4,-16,8,-11,-20,20,16,-2,-11,10,-19,-24,-6,-1,-18,-10,1,-7,9,-7,3,-22,-6,-18,9,3,19,4,-38,-18,-18,2,-15,-14,-10,1,-2,2,11,1,-17,-23,3,7,35,3,15,-12,15,-15,0,10,0,-33,-22,-1,-2,-22,23,-11,7,-23,-16,0,10,-1,2,-8,5,-12,25,0,-14,21,22,38,-10,-24,2,4,3,-20,-2,-29,-4,6,18,13,25,10,-25,-2,-5,22,-1,-41,9,-14,-6,-23,44,-5,-18,-6,-5,-38,-6,41,-3,-12,34,-6,-5,25,65,23,1,37,8,9,16,59,77,78,44,
24,38,11,11,22,19,10,-7,39,-2,16,7,17,14,6,26,-5,-13,2,9,-3,13,17,-9,8,33,9,24,-4,13,0,13,33,0,16,16,24,21,-6,17,15,6,-9,25,-2,1,-25,-6,13,-2,2,23,25,15,19,11,-18,-9,26,20,17,-6,32,5,-4,-4,2,5,38,12,22,-13,-29,6,10,20,2,8,0,23,-13,7,7,-34,-15,17,0,-11,6,5,9,6,29,23,0,-1,4,18,-11,-18,8,22,16,16,-22,10,-4,12,-2,16,25,13,-2,10,-11,-20,1,-3,14,10,-13,-18,0,13,3,5,9,19,-18,17,3,12,8,18,2,10,16,-20,12,11,16,13,5,-3,-7,1,9,19,19,22,47,43,23,-2,19,11,46,46,7,-28,15,25,36,13,-13,5,-27,-30,-1,-5,3,25,1,24,0,3,18,-7,10,23,14,-36,-7,8,2,12,24,-1,-8,18,15,11,9,18,16,-16,17,-19,-21,-59,-7,-17,-3,10,-28,-33,-49,-27,69,62,-33,-82,-85,-52,-60,20,3,4,-15,-8,10,-3,8,-28,19,30,36,40,-13,-14,-54,-9,20,9,20,-13,-24,-8,-3,-14,-43,-23,15,11,11,4,-6,14,12,26,33,46,-13,12,35,2,-8,-16,-9,11,6,-22,-30,-32,9,0,-17,3,-30,5,-12,22,-30,2,13,5,33,5,-4,-47,-32,-14,-2,10,-17,4,9,-21,10,-24,-1,-12,6,-9,-1,-5,-6,16,18,29,17,-19,-1,21,7,12,16,3,-30,3,4,3,-12,-8,-19,-10,3,6,24,-2,-2,-14,-22,-12,-26,3,-4,-3,-23,-26,-7,15,21,-15,-5,2,-17,20,3,-11,-26,4,-9,8,6,5,46,34,49,8,1,-5,13,61,72,49,27,-3,38,32,29,29,-30,-60,1,13,-10,35,9,-30,-69,9,-17,-33,4,-4,-17,-8,3,9,-1,36,20,0,-13,-8,18,14,45,28,18,27,
10,-12,-13,-15,-13,14,13,-6,6,2,-15,2,6,-9,5,4,-18,-18,1,8,-16,14,-13,-12,-11,7,-7,11,3,13,-8,-13,1,-1,-1,1,4,0,-8,0,-15,-1,-2,4,10,-14,-15,12,-14,-3,3,16,-4,11,-15,-17,-18,-15,4,10,8,-6,-12,-10,2,1,2,-8,-7,0,-18,3,-17,-9,12,-18,-10,-5,12,2,10,13,-9,-14,14,-14,7,6,-15,-10,9,-12,-10,-11,-16,15,1,-8,-9,11,2,-9,9,5,7,3,9,-5,-13,-15,-4,-9,-12,11,-10,-11,-13,-5,3,2,2,-6,8,11,0,-14,-10,12,6,-8,-2,3,-7,5,9,13,8,-14,9,-8,-7,-13,-4,3,5,11,8,11,-7,-3,-5,5,-1,-8,2,-14,9,-10,-14,-11,-8,-7,-16,-9,-13,-17,8,-12,-17,6,11,-17,-3,16,-1,-2,-3,-11,-14,14,-17,12,3,11,-12,-12,9,14,2,8,-18,-16,10,0,-1,11,14,9,-3,-10,-6,-10,-5,3,-6,6,-11,-15,-6,-17,16,-14,6,-3,-4,-5,6,-2,-3,6,1,12,0,-1,15,5,11,-16,16,-1,10,-1,5,-18,-6,2,13,-4,-17,12,-4,-3,-16,12,-13,2,13,-8,-2,14,12,-13,-17,1,-2,-1,6,5,-18,-1,-12,7,10,12,-8,3,-13,-12,9,3,3,0,-1,-19,-5,5,-5,-12,9,17,1,-12,-5,-1,0,-1,10,11,5,-14,15,4,-6,-2,12,-2,-6,-12,10,3,0,16,3,6,-4,-16,-16,14,-10,-18,-7,-12,0,-8,-8,9,-15,-6,-14,9,11,-17,16,15,1,-5,-17,15,6,-12,-2,-6,9,-10,-11,-11,-7,-14,-8,8,6,-11,1,6,-7,-7,-8,-11,7,-15,14,14,-13,-17,7,-16,-5,-9,0,14,10,-16,9,13,15,8,-2,-6,-4,-13,-5,15,-1,3,-7,-11,1,-13,-7,10,5,-11,0,13,-14,-6,-16,-15,15,-7,9,8,
1,13,14,-14,10,22,20,-17,17,9,2,-7,-6,26,8,15,-4,-7,11,15,8,-2,-16,-12,-12,-10,5,7,-15,-15,-5,6,25,24,-4,-9,-10,-11,18,-1,-22,17,7,-2,15,17,15,0,12,31,4,17,3,14,27,-1,-2,15,35,0,-33,-4,-42,14,34,16,34,35,32,-36,-6,-3,-32,-6,12,-9,-58,-7,-20,-33,21,30,-6,-63,-5,-19,9,1,-12,-16,-9,2,21,30,13,9,17,-12,-3,26,6,23,31,13,18,3,11,6,8,-4,-3,7,-14,-4,15,27,7,16,2,-9,-15,6,2,7,12,21,10,-23,-2,1,18,29,13,13,10,16,33,22,-11,2,21,-7,23,-8,-13,10,3,1,0,17,7,1,-19,-8,-11,-1,3,-3,-17,-37,-5,-4,-1,-4,-4,-23,15,-22,-3,18,-5,-23,5,55,-29,-2,-7,-24,1,23,16,-20,-8,3,-13,14,-27,-27,-10,-14,1,-7,-10,-20,-18,-14,20,15,17,-30,11,21,11,12,-7,-2,-7,15,0,-19,16,-21,4,10,22,10,-44,19,-12,-37,-5,39,-25,-77,5,38,29,11,-19,-55,-44,5,2,10,31,-6,-40,-36,13,-17,-9,-26,-38,-9,-17,15,14,-16,-15,-8,-9,-32,13,-2,10,-3,-50,-37,-78,11,32,6,28,-9,-9,-45,-4,-37,-42,-1,1,6,-70,8,-7,-22,1,34,-9,-55,-3,11,16,10,18,-38,-23,-7,4,-7,-13,-35,-48,-21,42,6,-7,-2,14,4,-3,0,-10,1,13,4,3,-4,15,8,7,27,-21,10,-15,8,-15,-10,9,19,26,6,3,-46,-49,0,7,4,-4,-7,-18,19,21,25,-39,-21,8,-3,13,22,-1,-5,-3,41,24,7,20,-10,-6,-62,12,3,-20,11,-27,-37,-75,5,4,23,17,-6,-40,-68,13,-4,17,-21,-13,2,-47,-1,-20,-61,-31,35,44,4,0,-26,-30,9,16,-2,16,-8,-12,27,-7,-6,-12,17,
9,12,23,6,-14,-9,-13,10,-4,16,20,-15,24,-24,7,15,6,24,4,-11,-6,23,15,25,-11,15,-2,6,-6,9,-17,-2,13,11,12,-3,19,-12,0,-6,-1,-6,14,7,-21,-18,13,-6,-4,22,2,20,-5,0,-33,-11,-11,-12,-15,-13,25,20,59,10,-21,-13,-20,-14,31,39,-11,1,12,19,-8,5,-13,-14,25,43,-24,-8,8,-21,-9,12,33,-10,-28,-22,-23,0,4,8,14,20,15,2,24,-13,-13,1,1,-13,-27,24,11,-14,-35,-22,9,-17,19,6,25,16,7,26,12,29,20,0,-6,-8,-22,17,-25,14,-10,12,-2,15,4,-8,4,-5,4,-19,-9,-32,12,-1,-3,18,-13,3,0,23,7,-1,24,5,-1,19,0,-1,32,-3,-21,-8,32,1,2,35,23,-5,-1,21,-1,15,35,38,-14,13,22,-4,31,10,14,19,1,-12,-6,1,12,30,16,14,25,21,1,6,27,14,2,7,7,-26,-43,-60,13,0,36,7,21,-29,-44,-23,59,45,11,-16,-4,17,29,48,44,20,20,-20,-1,-13,6,15,-13,-27,-46,-63,-13,6,-36,-11,-25,-37,-47,-50,-32,-43,7,-6,-26,2,-6,-19,-41,-14,-11,-5,0,11,-20,-23,14,-2,-24,0,23,19,43,-2,0,2,-18,-12,19,38,17,18,21,1,-14,19,-33,6,15,-18,-34,-6,-4,-20,-11,-20,11,3,-24,7,-25,9,-27,-25,15,-9,-38,-41,1,-16,-20,-30,-13,-22,-47,14,-6,-7,2,-13,-14,-11,2,4,-4,32,7,5,26,22,-22,24,-10,-17,-3,0,-16,-5,11,26,-8,-6,-40,-16,-5,11,7,-36,-37,-54,-7,10,3,-18,2,-2,-15,-7,-14,-17,8,20,1,-9,12,-23,23,24,39,53,30,-8,-5,-1,17,-4,-6,-3,-16,7,12,49,-29,10,-63,-17,23,28,45,-22,-4,-5,-26,6,44,18,22,0,4,-11,19,25,48,13,20,9,
-30,21,24,-1,-6,-6,23,0,1,-15,-6,24,21,21,22,-15,1,13,24,14,11,10,5,12,-11,0,-15,9,-9,-24,9,-33,-2,19,11,18,8,-16,-2,-7,-23,4,4,18,-19,3,-5,-16,1,1,12,25,4,-20,-12,-7,15,17,22,-12,-4,-18,-5,13,-8,-21,18,5,10,-65,20,17,6,21,20,18,-60,-9,24,7,-7,-4,17,-31,24,-10,-17,-22,-25,9,-16,27,-10,14,9,10,-28,-9,-17,2,10,-37,-16,-13,14,1,16,2,29,11,-7,-1,21,0,21,-11,17,23,2,-7,15,1,2,2,18,24,2,-2,20,-20,17,1,-15,-20,-32,-2,-2,-17,-16,-6,13,2,-11,2,-22,1,-28,-2,5,11,-4,20,5,-8,-12,13,4,-6,-20,-13,-28,15,9,4,18,6,31,-28,16,38,26,27,-4,30,-47,11,40,20,-11,29,5,-17,1,17,23,-15,-13,-11,-10,23,-5,5,15,-1,2,-23,23,1,-36,-17,-1,16,36,8,-24,-12,4,-15,-6,-8,-4,-17,-3,25,45,-11,-51,21,-48,-56,-34,-8,-26,-43,-25,-8,-37,-37,-24,-15,-40,-20,-17,-1,3,-20,-44,-2,15,-8,-5,22,-17,-25,-7,2,-1,-7,6,3,-7,-33,-7,16,33,18,13,-11,-52,1,17,-27,13,35,18,-62,22,19,23,-10,29,10,-72,8,19,0,-29,5,15,-57,13,-8,27,6,-13,-19,-22,36,1,0,26,-20,-13,-25,-9,22,1,-6,-13,-31,7,5,-8,3,13,1,-19,-4,33,12,27,-6,29,20,3,14,23,1,-12,26,16,2,-8,11,11,-17,28,21,-22,-8,4,-17,-7,-5,-33,-32,13,7,-2,-10,-8,-5,-42,-37,28,3,-11,-15,-23,-15,11,-1,12,-23,-25,-42,-14,26,20,25,1,8,28,-56,20,24,6,17,2,41,-62,6,39,36,16,36,26,-3,2,30,14,-6,14,-18,-20,9,-5,3,17,-2,-19,-8,
5,2,8,-17,8,-1,0,10,-16,2,19,29,-8,9,-5,-9,5,-10,7,14,10,1,24,-9,1,33,26,-2,7,-12,-9,-6,-9,-2,-9,2,-22,-6,-20,-15,-12,-1,8,5,7,-10,14,17,23,7,8,-4,-28,-11,4,14,5,-11,27,10,5,-12,7,-1,3,-32,4,-3,-16,50,1,7,-20,37,1,-30,11,-22,1,6,35,-26,-48,71,9,21,0,-18,-36,-7,-10,27,25,29,58,5,-7,9,-9,-12,-43,-49,-13,-15,-9,-8,-5,5,-14,0,1,-12,12,14,28,29,31,-4,-26,6,7,-7,-32,20,2,-22,-3,-3,14,-8,15,7,-17,4,-11,-19,-2,-4,-6,-11,-1,17,3,-2,13,12,21,6,-1,-31,-32,1,-11,3,-14,7,-3,-5,-4,25,16,0,12,-15,12,12,14,28,-12,14,-15,21,35,24,31,0,14,1,1,-18,-48,50,-8,23,8,17,3,-5,9,15,21,-4,22,45,42,5,-22,-17,-17,5,-44,-48,-41,-3,-3,33,42,36,7,-45,-16,34,31,54,18,-63,-23,14,3,28,22,-20,-61,-3,-19,10,29,3,15,36,29,-5,-18,-8,-22,-22,22,-24,-9,-13,-36,-34,-33,19,25,-31,-8,-11,-10,1,-4,-52,2,-17,15,-9,-6,4,-10,8,19,-21,-3,19,6,12,7,29,-4,41,44,-35,20,-10,-1,-6,-23,-47,-31,77,4,-6,6,-28,-19,5,-18,-4,-14,-27,-30,-2,-2,19,-25,-20,-38,-21,-19,-24,-36,-13,-10,1,-15,-3,-40,-23,28,-11,-1,8,33,1,-30,22,21,-3,-12,41,3,-1,-10,-9,7,28,-2,-13,-5,0,11,-2,12,-30,2,-7,1,14,39,-2,15,25,12,-37,-24,-24,-20,-9,-42,-15,12,-3,13,-43,-35,-20,-4,17,16,9,-8,-24,-3,46,0,18,-29,-13,59,6,73,-12,30,-18,49,43,-30,-5,-24,-5,33,12,-21,-28,-6,17,13,27,44,40,51,-7,
14,0,6,-4,-13,-31,2,-3,-5,-7,21,30,5,1,4,7,20,9,-4,6,-1,13,17,9,2,-27,3,18,-16,5,19,7,2,-25,-1,19,-22,5,-8,-16,2,10,1,-4,-7,18,16,7,26,-23,10,7,7,-27,-5,6,12,-2,-15,-12,32,0,58,-6,-5,-7,-22,-25,-22,23,-2,-6,29,-1,14,15,18,4,6,-11,1,-3,6,15,4,11,3,16,17,13,-5,-16,-30,3,7,25,10,27,-3,-3,-21,-12,-15,-12,12,-3,20,10,20,18,0,7,9,10,-1,7,5,17,16,12,-9,5,-9,-21,5,0,1,4,7,-4,-5,9,17,-5,-3,1,-14,-3,7,36,-14,-4,35,28,12,-13,14,7,12,-23,-8,-8,-23,4,-17,14,4,-8,-62,-2,25,-6,-20,-11,3,10,12,26,0,13,36,2,35,-2,36,13,6,10,-18,11,4,34,16,20,-15,-21,-3,30,8,-15,-17,19,12,-9,7,25,-35,3,-4,63,-11,-21,-48,-23,-5,9,81,39,16,11,-9,34,47,80,55,30,29,-12,21,55,-4,5,42,74,6,-21,-29,-28,-19,-1,0,22,32,10,4,-12,21,35,-14,19,38,48,16,9,17,-25,-1,20,14,4,-28,8,-18,14,-20,-16,26,22,89,-7,-1,16,-7,50,10,58,21,10,43,0,41,15,75,24,5,34,-24,0,14,31,7,7,13,25,-1,0,18,-14,20,13,37,15,22,15,-47,-25,-15,9,-20,-35,-12,-28,7,26,-13,38,8,4,19,0,0,0,4,24,25,15,-8,-5,-16,-8,-27,34,11,36,16,-12,6,-10,10,30,-4,5,19,18,30,39,-13,-24,6,29,30,2,14,-38,-28,-11,-37,-8,-31,21,-3,5,5,-20,-40,-13,42,21,-8,-13,-31,-43,37,74,13,-7,7,-39,35,22,58,32,9,22,-27,2,14,-9,24,15,-1,2,-19,39,-1,-8,-21,-23,-38,-21,25,-23,
-13,25,19,2,7,18,1,-13,15,-3,-2,-17,14,26,17,22,-10,9,-5,2,21,-1,-3,-6,4,24,1,22,4,-9,14,24,7,2,-15,8,-4,1,-14,8,-6,-9,2,-10,9,-15,7,15,-15,5,32,9,17,-3,18,16,5,2,41,6,-30,2,-21,14,18,-14,9,9,7,-7,18,20,20,25,-22,-10,-7,4,13,43,-17,9,5,68,-7,13,-1,-11,-4,-12,-9,-12,-15,22,-2,13,6,-10,21,35,40,8,1,21,34,-14,-26,-17,8,7,-9,-2,0,21,-23,10,-21,-7,-1,9,-4,-7,-11,-3,13,11,-23,-19,24,3,-2,5,-18,-28,-24,-13,-21,-7,-2,6,-13,-15,-8,-7,-9,20,-4,12,11,5,-2,48,34,-16,-6,-14,3,-6,9,-11,3,2,-5,2,0,28,42,-21,19,4,15,19,-11,33,-30,-24,26,23,-3,-13,-33,19,-8,5,34,-20,-8,37,-1,5,-14,13,11,14,14,9,26,32,12,7,22,20,37,-12,4,-26,-17,3,-2,-8,14,-38,-28,-18,13,-15,-49,-1,-20,-73,-54,-41,-10,-20,-23,-44,-28,13,-18,7,34,-11,-6,8,18,31,40,27,18,-11,-28,-12,20,18,-8,-4,10,4,16,6,24,-20,-10,-7,11,-1,-42,-22,-82,17,-14,-37,8,-10,12,-15,-10,26,25,22,-25,7,-22,-9,14,-2,8,-6,-20,62,-22,15,9,-4,-23,19,32,27,-6,3,-17,7,8,-7,4,2,21,22,-9,6,19,-25,1,-12,0,-21,-16,0,3,8,14,0,-32,13,-26,19,9,-14,20,13,13,16,-16,22,37,14,-26,1,2,-17,-1,-13,-11,-8,27,40,-12,-12,-1,-4,-10,-5,-25,15,27,17,17,12,24,-8,-24,-5,15,1,-29,-39,-53,19,23,11,6,0,-10,-12,23,24,-11,31,5,48,63,-23,35,18,22,-5,-9,42,-17,3,17,17,-47,-20,23,17,8,1,10,-7,-18,8,
1,-12,2,-6,4,31,17,14,-13,-12,-4,7,28,40,0,-17,5,13,11,-13,-24,19,15,4,-4,-11,-14,-16,-10,-11,4,-1,-3,22,-18,-26,9,-6,6,-7,0,-10,-11,1,-13,-6,-20,-20,-20,6,-13,-24,-3,-23,20,15,11,9,-33,36,0,-6,-33,-23,5,2,36,25,-11,-23,-6,32,4,16,9,11,46,-12,15,-23,-8,-11,13,17,6,15,6,15,-5,-12,15,8,22,1,0,-18,-16,-29,-4,-15,-2,9,-20,3,5,34,3,10,-4,5,-6,12,6,22,5,-1,16,-13,-14,6,18,-1,7,11,-5,-29,-4,5,10,11,28,15,-8,6,13,-13,-5,7,6,-25,-7,17,-10,-8,12,9,-35,-13,-38,5,-21,-56,-37,-7,0,-41,-13,43,76,79,-4,-7,-21,-8,49,70,43,-38,-17,2,-27,-1,-7,-34,-34,1,-11,-25,9,-20,-12,-19,-14,-15,8,16,7,-2,-3,-2,-1,-14,9,-1,-4,-31,-11,10,69,58,-2,-17,-32,22,79,95,22,-85,-128,-69,18,85,48,46,-55,-103,-43,7,-1,12,-18,-39,4,9,27,1,5,-13,32,51,47,-5,-22,-46,-13,-1,28,5,-2,15,-3,2,-9,7,-35,10,-17,4,-11,-48,-6,-13,46,0,-13,45,45,23,-67,-6,48,39,14,-10,-40,-28,4,20,4,12,1,-18,22,-11,-13,-7,-15,-26,19,32,13,9,-3,2,1,2,4,24,11,7,8,11,4,-25,8,-13,-15,9,2,5,9,64,-1,-11,3,11,-5,-5,22,-28,1,39,40,-21,-38,34,9,27,18,11,-4,-8,11,-1,21,1,1,19,-2,6,13,2,7,-8,6,-37,19,36,28,0,3,-29,-19,31,-36,-25,-16,-29,21,3,43,-24,-9,-10,5,28,9,-7,-10,-20,28,76,76,60,-5,6,11,32,41,4,75,14,-8,11,3,15,-9,-3,1,15,-3,-12,-2,-17,9,10,31,3,9,28,-31,-15,
16,2,-14,-14,-9,1,6,-12,-3,-11,5,6,14,12,-1,8,-10,4,15,-13,14,16,-16,-5,-17,-2,8,13,-2,-14,14,-12,-8,-3,-6,4,-13,5,-8,-15,-18,6,-13,-3,-1,9,10,-18,8,-16,10,-18,5,12,-12,13,15,-9,-6,-12,-15,-7,1,11,7,-16,-17,-12,-2,-9,-4,-9,-14,-7,0,14,-2,-4,11,17,1,2,-13,6,14,-1,-3,-10,10,5,0,9,-18,11,13,-6,13,-4,10,5,-14,-7,4,-10,1,10,12,-3,5,-13,-7,-1,10,-13,3,1,-1,12,-14,-17,-8,-19,0,6,-8,-1,-1,9,-11,16,14,-9,13,-17,15,16,-13,-15,-7,-11,7,12,-3,-1,13,14,-17,-4,14,-4,-12,1,-7,6,1,-17,-13,-11,-15,-8,-8,10,-16,-13,10,-6,-12,16,-11,16,2,-13,6,11,-6,-8,-17,-6,14,-9,-2,0,15,-16,1,-11,-14,-16,-8,12,2,6,-17,-14,5,-16,-9,16,-6,9,5,-11,13,-16,7,-16,5,-15,-17,11,8,7,5,-14,7,-12,13,9,8,10,-8,4,-18,3,-8,-13,15,1,3,-17,-16,0,-5,-13,2,-11,7,-6,14,14,11,-4,10,13,4,-8,8,13,15,2,-8,-13,-16,7,0,8,-4,8,12,-14,6,14,-5,11,-10,-14,12,-11,4,-3,-12,16,3,2,13,-7,-9,13,-3,8,6,-5,15,0,-4,-7,-2,-9,-7,6,4,15,12,1,-3,-6,-3,3,-2,-7,-6,-4,8,3,0,6,-15,0,1,11,0,-14,8,-2,-19,-10,-5,-6,-13,3,-2,-10,11,-17,13,-5,-6,-3,8,16,-13,1,5,-14,-1,2,-11,-3,-14,15,6,9,-15,11,-15,8,1,-3,-11,6,-16,-8,-6,-17,5,-15,-10,11,-3,6,0,-16,-4,-10,2,-5,-3,-11,-19,2,-3,-2,-13,2,11,2,15,-18,5,-17,-9,-5,15,-12,-6,-2,-1,-10,10,10,-1,-4,
16,27,-8,-6,-2,-9,13,-2,24,-5,-1,-10,-13,20,6,14,-1,19,5,17,-8,-28,-14,8,31,25,-27,-20,11,-47,11,-6,-6,-6,-17,-15,-22,5,14,15,5,-14,2,-6,-12,12,12,-9,1,-14,29,19,16,-11,-19,31,29,14,9,-5,-17,17,0,4,-1,-16,13,10,-14,3,-11,-39,-5,23,-8,-28,8,-31,-2,15,-7,-20,-28,2,-41,-21,15,-9,10,4,-33,-7,-12,-15,-29,-8,11,16,3,9,17,-2,3,10,-10,11,1,-2,-10,-12,-9,23,9,-8,-12,-14,5,23,0,-23,6,6,4,-6,-18,-32,-33,-50,1,11,-9,-3,-50,-20,-26,-11,10,-1,7,-8,-12,-47,-27,-6,16,5,-3,1,2,-5,-7,-6,14,-2,21,11,5,23,20,20,-9,-9,14,-17,8,2,-10,-12,-17,-6,28,29,8,-27,15,-22,-11,26,-12,-18,-31,5,-7,-10,28,-8,8,17,21,-11,-24,-4,34,-2,13,20,12,26,10,9,15,24,38,-4,6,-11,-22,-35,5,4,16,24,-13,-41,-14,5,20,4,-16,12,15,10,10,-14,-38,-37,-23,-26,4,-11,-19,-54,-46,-7,21,-2,0,-38,-12,-48,-10,2,24,20,12,-6,21,2,21,-11,8,-8,14,1,1,8,14,-16,-25,-15,-1,-18,26,7,-24,-4,-19,-28,9,7,15,-25,14,-51,-14,14,18,10,-25,3,-53,-44,24,19,-2,-4,-22,-23,-47,1,21,24,22,25,-11,24,5,16,-9,9,-7,5,27,17,-4,12,-2,9,8,0,11,12,21,-7,-1,-22,-1,-9,10,-1,-34,-30,-15,-53,-4,10,4,-24,-28,-60,-42,5,-15,9,-19,-6,-44,-46,-33,10,3,20,-6,-3,32,-7,9,0,24,-11,-12,-3,-16,-4,6,21,14,-1,-15,3,14,23,-7,-13,-17,-33,9,10,20,-28,24,-41,-40,24,9,-16,-33,-2,-61,-6,11,-31,-18,-13,-6,-28,-49,-2,8,-13,-13,-21,
0,-17,-11,-3,11,6,12,-4,16,0,-16,-2,16,-2,8,-16,-14,14,0,-10,-27,0,6,8,4,13,14,9,-1,-12,-23,5,0,24,-9,-15,-13,-8,-2,13,-23,-9,-6,19,0,-13,-11,-31,-9,4,-24,-22,-9,-11,3,-6,22,-10,-23,-2,49,5,4,4,0,-1,39,17,10,-15,-9,20,-1,2,27,52,8,-21,-26,-26,3,-3,4,-58,-9,-21,18,7,-2,-1,10,19,39,14,12,-10,-23,6,5,-16,-10,-10,-9,4,-17,6,29,6,-16,1,2,11,-4,-7,30,-13,15,-5,-14,18,-3,27,-8,-7,22,-14,17,23,0,17,46,46,-14,-9,11,-9,18,-10,-12,-37,-6,11,-3,10,-3,-12,-36,2,-12,-17,9,-43,-17,-27,16,6,-7,24,52,52,-26,-4,0,21,18,-7,-15,-2,-18,3,5,-5,-3,-26,-23,1,-4,6,20,21,15,-7,14,-17,-6,20,20,-47,-24,-5,-1,4,6,-19,-16,-17,-24,-38,4,-45,-36,-28,-31,25,48,80,5,-42,-68,6,20,21,19,1,-44,5,8,0,44,22,21,22,25,-6,13,43,15,24,43,20,-25,-18,-10,-30,-30,-24,-48,-51,9,10,0,-8,-30,-27,-20,3,-15,-8,-15,2,-16,26,13,15,-8,23,46,47,12,24,33,31,19,3,-53,-20,-5,6,-1,6,26,-1,-21,0,5,-10,-11,28,15,-59,9,5,1,24,21,-18,-20,9,-6,-5,-13,-27,-30,-52,11,-1,-22,-4,-11,12,-1,36,25,-17,-27,13,9,17,40,-3,13,29,42,-5,-45,13,17,31,16,27,25,-5,-11,7,5,11,30,4,-10,-15,2,-4,28,-18,-24,-72,7,15,19,26,-1,-19,-15,7,-24,-29,16,3,-19,25,14,-1,-2,-4,49,45,34,5,-15,-18,12,53,19,-13,2,-12,26,14,9,-16,-47,-14,-31,-5,20,8,13,-11,5,0,8,-8,42,-8,-18,13,12,20,51,38,9,-23,
12,3,-8,7,5,18,11,3,0,-8,-8,-18,0,8,21,0,10,20,-1,32,22,17,17,26,-13,12,1,20,3,-10,0,20,-13,-14,5,9,-12,-5,10,12,-8,-12,4,-10,-27,2,16,-10,-17,1,-13,2,-3,-12,12,1,-5,-3,-22,2,-12,6,-45,-10,42,28,22,6,-21,-29,30,30,33,-9,5,-20,1,-2,13,36,-5,26,-4,30,-6,14,22,3,-12,-4,-7,-16,-36,-8,-20,-10,0,6,20,37,23,-10,12,-1,28,15,1,-7,-3,-21,-14,-6,-18,-14,2,4,15,1,-14,-4,25,19,15,-5,16,-2,-5,1,23,8,-9,15,19,-8,-31,1,-5,11,-8,-1,20,-25,-17,-12,16,-4,-2,17,-16,-1,16,25,13,2,8,-2,15,26,20,28,-15,14,13,-2,28,13,15,-9,29,30,2,4,6,0,-15,17,21,29,-20,-15,14,19,-17,1,31,-11,-6,0,-6,-1,-3,24,-4,-10,-11,16,21,53,6,25,33,33,17,-31,-27,-89,-46,-10,-6,-21,-7,-7,-62,-10,-19,-25,-49,13,-16,-52,-44,-22,5,-43,-23,-22,-24,-51,-9,48,34,1,-13,3,4,10,27,-12,18,-8,20,-8,14,8,-29,-14,-20,10,9,7,-4,-19,-3,8,-13,-4,-40,-3,-80,-25,26,1,-46,-48,-36,-28,16,29,-13,-19,8,-7,-32,-8,-5,-4,-49,-11,17,43,-4,22,10,7,0,0,16,6,-12,24,-13,9,-15,-18,7,-8,11,15,13,10,20,2,-32,-12,24,-6,-32,-37,-5,10,9,14,-19,23,6,-6,45,30,0,-16,4,20,23,0,18,-2,10,10,9,20,-27,15,5,16,12,-13,19,-28,-17,-36,-14,-57,-10,-18,-12,14,31,17,32,-25,-30,-8,21,49,22,19,-79,-13,4,14,56,32,1,-30,6,32,30,22,-2,24,32,-9,26,71,13,-19,15,27,-11,10,6,-23,-34,-16,27,18,-20,-27,-46,-93,-54,19,
34,-10,16,18,-7,3,1,-6,-5,0,2,13,11,-10,-18,-14,-4,0,1,-9,-16,-6,-5,-16,-13,-22,-10,-11,3,-3,7,23,7,-17,-4,19,18,4,15,15,-4,10,5,-14,12,8,7,24,18,36,9,-2,-19,-17,5,33,1,6,-20,3,10,7,17,4,-9,40,5,-21,-17,-3,-7,-13,19,-12,-12,-17,13,28,-30,-16,22,9,17,5,-3,-10,5,21,37,31,27,4,0,-21,-35,3,26,34,16,0,18,38,28,20,8,9,3,-9,6,18,7,-17,0,-10,-3,-6,8,5,18,-18,-6,16,17,-16,-7,-7,24,-1,10,-7,-1,-25,11,4,28,25,16,38,2,27,9,-16,24,8,30,20,32,23,6,-4,-3,14,18,15,20,0,1,24,1,17,28,-3,8,23,12,-5,-26,41,23,-6,18,-9,-3,-3,58,2,-33,10,-2,17,9,23,0,-8,-13,8,-12,3,27,-14,14,-1,-17,-6,9,11,-13,36,63,49,31,7,2,-17,-30,-36,-17,18,-8,2,-10,-7,-20,-9,23,37,36,-3,7,34,27,22,0,15,27,24,44,11,-4,-37,-43,36,29,45,20,13,8,22,-8,17,39,29,30,32,31,5,4,4,-23,6,25,11,6,18,-2,-14,8,-4,34,9,-1,34,7,-5,-13,31,0,-15,-8,-14,-3,-29,29,8,-28,3,33,-1,17,-37,23,17,8,11,34,-3,-4,-20,-3,21,12,-4,2,11,24,-9,5,-3,0,-11,-6,-1,6,-5,6,-8,2,1,-26,-13,14,7,-1,-18,-9,-20,-22,16,0,-29,-19,10,-5,-29,-32,9,9,-15,12,16,13,28,26,24,32,25,-13,4,-2,31,8,4,6,41,-18,17,6,13,-10,-24,-6,-4,-11,20,25,8,-1,-18,-8,0,12,-14,-53,5,-7,-15,15,-27,-14,-32,34,22,-38,-8,-9,1,22,7,11,-3,-20,-2,7,26,48,0,-1,12,-54,-27,8,36
    );

    constant FC1_B_INT: integer_vector(0 to FC1_N-1) := (
-16,-19,11,16,3,-12,-6,8,13,6,-8,17,-13,-15,8,3,13,28,9,-18,-15,-5,-24,33,22,-12,-13,4,-2,-3,1,2
    );

constant FC1_W: mem_t(0 to FC1_M-1)(FC1_N*FC1_DTW-1 downto 0);
constant FC1_B: mem_t(0 to FC1_N/FC1_P-1)(FC1_P*FC1_DTW-1 downto 0);

end package;

package body fc1_rom is
    -- with change ColRow
    function intv_to_mem(intv: integer_vector; constant DTW,P,M: positive) return mem_t is
        variable slv: std_logic_vector(P*DTW-1 downto 0);
        variable ret: mem_t(0 to intv'length/P-1)(P*DTW-1 downto 0);
    begin
        for i in ret'range loop
            for pp in 0 to P-1 loop
                slv((pp+1)*DTW-1 downto pp*DTW) := std_logic_vector(to_signed(intv(M*pp+i), DTW));
            end loop;
            ret(i) := slv;
        end loop;
        return ret;
    end function;

    constant FC1_W: mem_t(0 to FC1_M-1)(FC1_N*FC1_DTW-1 downto 0) := intv_to_mem(FC1_W_INT, FC1_DTW, FC1_N, FC1_M);
    constant FC1_B: mem_t(0 to FC1_N/FC1_P-1)(FC1_P*FC1_DTW-1 downto 0) := intv_to_mem(FC1_B_INT, FC1_DTW, FC1_P, 1);

end package body;
