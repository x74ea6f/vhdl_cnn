
library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.piping_pkg.all;

package fc1_rom is
    constant FC1_M: positive := 8*7*7;
    constant FC1_N: positive := 32;
    constant FC1_DTW: positive := 8;
    constant FC1_P: positive := 1;
    -- constant FC1_P: positive := 4;

    -- function intv_to_mem(intv: integer_vector; constant DTW: positive; constant P: positive) return mem_t;

    constant FC1_W_INT: integer_vector(0 to FC1_M*FC1_N-1) := (
5,4,6,-1,-1,-2,4,-7,-6,2,8,6,-8,-5,-2,4,0,8,8,9,0,8,12,-1,-2,-1,10,8,-12,4,13,-5,-1,-2,9,-1,0,7,3,-9,0,8,-8,0,0,1,-4,-3,-2,6,4,7,5,12,7,-3,-3,2,8,11,4,-1,3,4,3,3,22,9,-24,-6,4,4,6,-3,-2,-8,3,-1,-6,-5,4,-1,3,3,6,-6,-2,3,-3,9,2,4,3,7,5,3,2,5,2,3,8,4,-7,-11,-5,-8,-9,-1,2,12,-6,-14,3,4,1,4,-8,7,9,0,-2,5,-5,-10,-1,11,-5,-8,3,4,-2,1,10,3,-4,-3,4,-5,5,3,0,-14,-13,-11,-4,0,-1,-4,3,1,-6,3,5,3,2,-12,-16,2,16,6,-2,4,3,1,23,15,16,-21,-3,-2,0,0,-8,1,-5,5,5,3,-8,-10,-6,18,7,-3,4,2,1,14,8,3,8,10,-3,4,-7,-1,0,-1,-2,0,3,-2,-2,-1,1,4,14,7,7,-3,10,11,9,11,-2,0,1,-7,0,22,-4,-16,-28,-9,-8,-12,-18,-14,2,4,-1,-8,-40,-19,0,6,19,9,0,-1,-5,2,7,1,-5,-4,-15,-2,-3,6,-4,-11,0,-10,-1,-2,3,4,-12,-5,4,-2,0,-20,3,6,2,7,-4,-6,-5,-2,6,5,10,22,9,8,3,10,-1,8,7,-10,-7,-1,9,1,-5,0,-8,-9,-4,-11,6,3,-5,4,-3,-5,-3,0,-3,-21,-7,-2,-2,8,2,-11,-2,0,5,8,3,-1,-13,-21,-6,-12,8,-12,6,8,-9,-5,-12,4,-3,7,9,26,-1,-2,-6,-11,6,-1,-2,-11,-1,9,-7,7,7,6,11,11,1,4,-5,-6,-8,12,9,-4,-24,-5,-3,12,19,14,3,-10,-1,6,-5,-15,-9,9,21,-1,-5,-9,-17,-5,3,9,3,7,1,-3,0,10,16,-25,-1,1,-10,2,6,7,
-1,4,-5,-5,-6,-3,4,-4,-1,11,4,-2,-6,5,3,6,4,-5,-3,0,9,-5,2,-5,-15,6,3,4,-10,-6,-5,3,-4,3,-11,4,3,14,8,5,10,-2,0,6,-1,5,8,0,8,7,-3,3,-1,10,8,3,1,-1,-9,4,5,3,4,6,9,-1,-4,-6,-15,5,0,4,14,9,-8,-6,3,4,-23,-17,-5,-2,10,11,1,2,-11,3,-1,4,6,6,1,2,4,12,5,2,0,1,4,-4,-8,3,4,1,7,8,6,-6,-2,3,8,-4,9,6,-1,-3,-2,-7,-10,-12,-5,-2,3,8,-1,-9,-7,1,-6,-4,0,10,1,2,6,13,15,0,0,-20,-9,-3,0,-1,6,3,4,-7,-9,0,9,-5,1,-3,-3,-5,11,11,-9,2,10,5,-1,-4,-1,-7,-2,1,-2,9,5,-6,1,-8,-8,-20,-17,-8,-8,18,4,-2,-2,3,1,17,5,11,11,11,0,8,11,5,4,1,9,4,3,4,2,9,9,-2,7,-4,-3,-4,-1,-7,-13,-14,-4,-3,1,-1,-4,0,2,-33,-27,7,-1,-10,-7,11,-7,3,4,-7,-5,-2,16,22,31,18,7,-7,-22,-6,6,7,-3,0,-11,8,-3,-3,-1,5,3,9,0,-2,-2,-6,3,3,12,1,0,0,2,8,-4,-2,-8,-6,6,7,-5,8,-2,6,6,6,-5,0,4,3,11,10,2,-4,4,3,5,6,-2,1,0,11,-3,8,5,2,-4,-2,8,-3,5,-6,25,10,1,2,5,-3,2,27,15,5,5,5,5,-14,8,-12,5,-3,-1,6,-1,10,-12,-1,0,3,8,14,5,-3,6,8,6,0,-12,-8,-11,-5,1,0,3,-4,-5,2,1,6,3,11,1,12,-2,8,1,10,-2,8,2,-7,-10,-2,-2,-6,-1,-6,-4,2,8,-11,-11,-16,-13,-6,-11,-4,3,7,11,11,11,12,-6,-11,-6,11,9,8,15,19,
7,6,2,-6,-2,3,2,-3,-1,2,-5,1,-3,-3,-10,-4,-3,4,-4,-4,3,-2,11,5,6,4,-9,0,-9,4,7,9,-2,5,4,-2,-4,-3,4,-3,10,2,-4,5,-2,-1,-3,5,-6,8,8,1,7,0,5,10,0,3,-20,0,6,16,6,-2,1,-3,3,13,18,0,0,6,-8,-6,1,-1,2,8,-3,-4,-8,4,2,-1,8,-10,-6,-4,6,4,0,13,5,2,9,4,0,7,4,6,-3,-2,-4,0,0,-7,0,-2,-4,-1,2,-6,-7,6,7,7,1,-5,2,11,8,-7,-11,2,-6,-2,1,-4,-9,-2,1,2,0,6,7,-5,6,-5,0,2,-17,-19,-11,-9,6,0,5,4,0,-3,-3,17,5,1,-3,14,10,-8,-15,-10,1,-11,1,0,5,-3,8,9,-3,0,-6,-1,0,-3,-4,-2,-4,3,-4,-2,0,6,8,0,2,1,5,9,0,11,11,10,9,5,1,1,-2,0,-2,3,1,2,8,-4,-1,-2,-7,6,9,-2,-2,-4,-10,11,11,9,14,1,17,19,8,10,2,-3,12,-2,-18,-26,8,11,0,6,-7,-23,2,8,1,-3,0,0,-7,0,6,-2,3,1,3,5,1,5,-2,-2,8,4,4,5,1,-3,2,0,1,8,1,-2,-2,-7,2,0,8,1,-8,-7,-3,5,6,16,15,-3,0,4,2,9,9,-1,1,-1,-3,5,-2,-5,-11,-1,0,7,8,5,1,15,-1,-9,1,-2,11,11,6,-6,8,-4,4,7,35,28,10,-9,-4,1,-11,-4,24,8,2,-12,6,-9,7,16,5,-2,3,2,-1,42,16,7,5,0,-4,5,1,2,-1,1,4,5,9,3,-1,9,8,9,-4,10,7,-7,1,-6,3,-3,2,0,11,2,1,4,9,3,-13,-13,-4,-4,10,-3,-11,-9,-8,1,3,7,7,5,-3,-2,-2,10,4,-17,3,9,1,8,9,-3,
-7,-3,-1,-3,2,3,0,-2,-4,-7,4,3,5,-1,3,-4,0,3,0,1,5,2,5,-3,-5,2,-5,5,1,-4,-1,2,-5,1,2,3,-4,-5,-1,-4,1,-4,4,-1,5,-5,-5,-5,-2,5,5,-2,2,0,-1,1,-3,-2,-5,3,2,6,-5,-6,1,2,-3,0,-2,5,-6,1,1,3,-4,2,-6,-1,-6,3,-5,-3,-1,-2,-6,-4,-3,-4,0,-3,-5,6,4,5,-4,0,-1,-2,5,-5,-3,1,-6,-1,1,1,-6,1,0,3,0,6,-5,-3,-2,-7,-2,3,-4,5,1,-6,-3,-2,0,6,0,5,-4,0,3,-4,-7,-4,1,-5,3,-3,5,4,0,-5,6,-2,-5,-3,4,0,-4,1,-7,1,-3,1,-1,-6,-2,-5,5,1,-3,-6,4,1,-4,-6,-2,-2,-7,-6,2,-4,-6,-2,-3,-3,2,-3,2,3,6,-2,-3,6,-7,-3,5,-2,4,3,3,-6,-6,-5,3,-4,6,5,3,0,3,4,0,-3,-1,-2,-1,-1,-2,6,1,4,-2,5,-2,-2,3,3,-5,-3,-3,-6,2,4,-5,-5,0,0,-6,-1,-3,3,-6,3,-1,-5,0,-7,-2,-4,-6,1,-6,-2,-4,5,4,-5,-6,3,6,6,4,-5,-3,-3,6,-5,6,-2,-6,-2,6,-1,3,3,-2,2,-3,1,2,0,-5,-2,0,-4,1,-4,-6,-3,4,0,-3,5,2,-5,-6,-6,4,-2,-1,-4,2,-6,3,-1,-3,3,0,-6,-3,-2,-1,-5,-2,-3,0,-6,4,5,-3,6,-2,4,-6,6,3,-3,1,5,0,5,5,1,-6,0,-2,-7,1,-6,-4,-5,6,-2,-2,5,-6,2,0,3,3,0,-6,-2,3,-2,-5,0,2,1,4,-7,-1,4,2,-1,-5,5,4,-5,6,-5,5,1,2,-6,0,4,-1,-3,-2,5,6,0,-7,3,3,1,5,-4,-2,-3,-1,-1,-7,3,5,-4,-5,2,3,2,
5,2,-3,-5,2,1,-7,-2,2,1,4,-5,-3,-1,-1,-5,-4,4,-3,-3,1,-1,-5,3,5,4,5,4,-5,2,-4,3,0,-4,5,5,-4,-7,1,2,2,4,0,-2,-3,-1,-7,-1,-6,-3,4,2,-4,-4,4,-4,0,-7,3,-4,5,-3,-5,3,2,-6,-5,-6,0,-2,-4,5,-5,-1,0,-1,-7,-3,4,2,-1,-4,-5,-4,0,5,5,-2,-6,5,-7,-3,-3,4,5,-6,-5,2,-7,3,5,-7,-1,5,2,5,-8,1,0,-7,-5,-6,-1,-2,1,0,2,0,3,-7,-7,0,-6,5,-2,-6,-2,-4,2,0,3,0,-1,-3,-6,-6,-5,-5,-4,-4,-5,5,-4,-1,-7,5,0,2,2,5,2,0,0,-5,-4,-7,-5,3,-4,2,3,-3,2,2,5,2,-5,-2,1,-6,0,5,-5,0,4,-1,-4,-2,-2,-1,2,-6,3,3,-5,-4,4,-4,-8,-2,5,1,3,-4,5,4,1,-1,3,2,-2,5,1,5,-2,0,3,-3,3,2,-2,-7,-1,2,-1,4,-3,0,-4,4,-2,-2,2,-6,-2,-4,-3,2,-3,2,4,-5,0,1,-3,6,-2,2,-7,0,1,-6,1,5,0,-6,5,2,-6,-4,-6,5,1,4,-8,3,-6,-6,-5,-1,4,-6,4,-4,2,-6,4,0,-4,-3,3,-4,5,2,5,4,-5,-4,2,-6,-2,-6,-4,-4,0,5,-2,-2,-6,4,2,2,-6,-3,0,4,-1,1,-1,-1,0,-4,1,4,-2,0,2,-2,-4,0,6,-6,-4,-6,-3,-2,1,4,6,5,-6,-5,-3,-3,6,-2,-4,5,4,5,2,-6,-6,4,-6,-7,-3,0,6,3,0,-5,5,-6,2,2,-4,5,-2,1,-4,-4,2,4,-2,-2,-3,-1,0,5,3,0,0,-6,-2,-3,-5,1,1,3,-2,-4,1,3,-7,-7,2,-1,5,-4,-1,-8,-6,3,2,5,5,-1,-4,1,-6,4,
-3,1,3,-4,1,-2,2,9,22,17,1,6,1,-2,22,12,3,9,0,0,-12,12,-8,0,4,-11,2,-19,7,-2,-10,-11,-7,11,-7,6,11,3,-1,-1,5,4,6,1,13,9,2,4,-5,-10,-8,-15,1,-7,-13,-3,-6,-4,8,9,2,-1,-5,2,10,26,24,13,11,8,-4,17,9,0,5,-8,-8,-15,10,17,-5,1,-11,-12,-12,3,-7,-8,6,0,-14,-7,-4,-5,2,-4,-5,-9,4,5,4,-1,-5,0,-4,-6,11,24,13,15,9,5,5,5,-2,9,9,-5,-10,-2,-6,-8,5,2,4,-19,6,5,-3,-11,-5,8,-9,-3,2,13,-6,2,-10,-4,-8,13,12,13,1,-4,-3,1,-5,2,-3,-14,-14,-4,3,9,17,5,-2,-1,2,2,12,8,14,16,2,16,-2,-7,-5,-6,11,5,-8,-2,-8,-1,-4,12,6,-22,7,-1,-13,-6,2,-5,-8,-1,3,2,6,-1,-3,-4,-6,-2,-5,-5,-7,0,-10,-5,2,12,12,10,0,2,-2,-12,3,11,7,-7,-2,-1,10,7,5,23,33,8,3,33,15,25,-8,-15,-3,-8,21,24,11,-10,-12,-5,-10,-5,-9,0,-10,-11,-7,-3,12,11,-5,-6,-3,-8,-6,14,13,6,4,7,3,5,6,-4,7,6,-8,-19,-1,-22,-18,3,-2,9,-6,-8,-7,-7,-14,-1,12,0,1,-2,1,4,5,3,-2,-9,4,3,16,2,-4,-3,-7,-3,-5,-16,-11,5,-11,-3,-8,-25,-18,-13,-4,-10,-7,-1,-38,-29,-19,1,-9,2,1,-31,2,-5,5,-1,-2,11,-38,-8,-7,1,-5,-6,4,-47,-29,2,-13,-7,-8,-4,-10,-8,6,-4,2,-10,-7,-7,-11,-3,-5,-11,18,21,16,8,9,-6,1,17,11,16,25,19,3,13,-9,-12,-2,3,10,-13,-24,6,-3,2,3,6,8,-10,10,-1,-4,-10,-9,-10,-9,26,15,16,2,1,-3,-11,
0,2,12,-1,11,9,2,0,4,2,12,11,-3,-2,-2,9,-3,0,5,4,0,-4,-1,0,11,2,8,4,5,-6,12,5,-7,6,1,3,-1,6,8,12,10,-7,1,2,3,-5,5,6,-9,-6,-4,2,0,1,0,4,7,10,4,-11,5,-8,-2,-3,-2,-2,-4,-2,-6,-1,3,-5,-13,-4,15,9,-8,-4,-14,-5,8,2,3,1,-5,5,7,12,0,4,-1,1,-2,6,11,3,-4,3,3,4,-6,4,13,0,0,-4,3,-5,10,4,-5,-11,-1,-4,-12,-8,1,-1,5,8,2,3,19,8,3,1,-9,-5,2,3,2,-3,-2,-1,5,14,15,12,2,-4,3,11,3,-5,-7,4,6,-3,5,16,5,13,5,1,0,-5,-13,-4,5,4,-6,-3,-5,-5,-6,-7,1,-17,6,2,0,4,-2,11,-7,0,9,4,16,15,5,-3,-6,0,10,4,5,0,-1,-6,-6,11,4,12,0,-1,4,-1,1,1,-1,5,-5,-4,-6,-7,-6,0,-1,-4,0,0,8,-8,-3,7,-6,-5,-10,-9,-4,15,3,-7,-9,-12,-21,-6,3,-14,-5,-5,-5,-5,22,-10,-6,7,7,-1,20,15,5,-8,-6,-2,22,9,13,19,10,-2,-5,-8,-10,5,-10,-8,-8,-2,0,4,-1,-5,5,8,-1,13,8,20,6,5,11,2,-1,2,0,-4,9,7,3,4,5,-10,6,-4,-5,-6,-3,-3,-5,-4,0,-14,-2,-1,2,3,3,0,8,3,1,-4,-5,6,2,1,3,-17,-22,-29,-19,-4,7,2,15,4,-23,-14,-3,6,-4,2,7,-6,1,-6,4,6,4,-11,-18,-11,-1,-6,1,0,-29,-21,-4,-6,7,3,2,15,7,2,-3,-7,5,-10,-7,9,9,10,-1,0,-9,-13,-17,-14,-5,-18,-1,1,3,5,21,9,0,-3,6,15,5,8,5,4,6,3,10,15,20,10,-6,1,0,-1,-8,-1,9,-3,
2,-2,-7,-1,-2,-3,10,11,1,6,7,1,6,2,-2,0,7,-8,-9,6,10,11,12,12,1,19,13,-5,1,7,6,4,18,2,-6,1,-7,-7,-11,-4,-11,-4,5,2,3,4,10,-5,-6,-3,6,-2,-4,4,1,4,1,8,11,6,-11,5,7,-1,-1,-6,1,-17,-7,5,7,4,14,-2,-2,4,0,8,0,6,10,15,11,0,-3,-4,-8,-5,-10,0,3,3,-3,-8,-5,4,-3,8,-4,3,5,12,3,-3,5,1,-4,9,1,1,5,13,-3,6,12,9,-7,9,2,-2,5,7,8,5,16,-2,2,5,-4,5,2,-9,-2,1,-3,-14,-12,0,-3,2,-1,-3,-1,12,14,5,-4,-2,-8,-8,3,1,0,-2,3,6,13,10,18,17,7,-3,2,9,-3,8,-9,-7,-1,4,12,9,-1,3,1,-2,8,3,12,19,5,0,0,-4,-6,-7,-2,-8,-4,1,-6,-3,6,-3,-5,2,1,2,4,4,1,-4,-2,-1,-3,8,10,5,5,1,-3,5,-9,-2,-20,-10,0,-1,-2,6,-3,-26,-7,-2,-4,0,3,-2,-17,5,6,6,-16,-24,-33,-13,-5,4,10,-1,-7,-32,-1,4,1,-4,-3,-18,-3,-11,-9,10,2,2,9,6,3,5,1,1,9,22,6,9,16,-6,6,5,10,12,16,5,-15,-1,7,-2,0,4,-17,-18,7,3,-9,0,-2,0,-9,8,-2,-3,2,2,0,-10,-2,-3,0,7,7,5,-4,-1,-2,6,-4,14,3,6,-3,15,22,3,-6,4,5,4,-7,22,-17,0,-7,4,8,-9,14,-4,2,3,4,5,-10,16,21,10,-2,9,6,6,18,17,12,-1,-4,7,2,-6,-7,0,5,-1,5,-4,6,8,4,-7,5,5,12,13,-5,-2,-1,-9,8,12,3,8,8,9,-5,-7,-5,11,13,7,11,-17,-5,-9,-12,-3,-13,-10,-17,-6,-3,-1,2,4,4,-1,
13,6,-12,-4,-14,-11,3,13,0,-8,-10,-2,3,7,9,-6,8,4,16,10,-1,-8,13,14,3,6,8,-5,5,9,3,-5,8,8,-3,2,3,2,3,-1,-7,-13,10,1,-3,-2,-4,-2,-8,12,13,9,5,10,9,6,7,9,0,-7,-22,-17,5,8,18,-3,-12,-22,-14,0,12,-9,1,3,-12,2,6,11,14,13,-2,5,12,4,11,3,-3,2,4,-3,8,2,3,0,3,0,10,2,12,2,-1,1,-5,1,-6,10,6,4,-7,4,3,8,10,-1,2,0,10,8,-2,4,6,15,-6,-1,12,6,-6,1,4,-2,5,1,1,5,-2,-8,-4,3,0,-3,19,15,4,5,1,7,7,7,-6,-2,3,-1,2,10,8,4,4,4,11,-6,-8,12,-4,-4,7,5,-12,-15,7,10,-1,7,10,-3,-6,11,2,8,2,-7,-4,-6,-1,3,-4,-3,-5,1,1,10,-2,2,3,-4,0,0,3,11,11,-1,5,12,4,11,14,-2,6,9,7,9,6,12,18,2,-21,-19,-2,2,-7,-14,-26,-36,-24,0,-8,-9,12,14,-17,-7,-3,14,21,27,-10,11,2,9,5,9,-5,-6,6,15,5,9,-10,-13,-7,-10,-3,-9,9,-3,-8,2,11,7,5,15,2,-6,7,14,18,-2,17,8,12,7,10,1,1,5,1,-8,-7,16,-1,-13,7,2,-3,15,-7,7,-7,7,5,21,0,1,7,1,5,0,2,7,5,4,-3,-4,5,10,28,23,1,17,5,6,8,9,33,14,11,5,2,13,0,7,8,3,-4,15,30,17,-5,2,5,-4,-6,6,17,1,8,6,1,4,42,30,12,4,-2,9,-2,2,-2,4,3,13,4,-8,2,0,-13,-12,-9,9,-3,-13,6,-5,-6,-14,0,5,0,-6,-9,-7,-6,7,9,-1,-8,-6,10,1,4,-13,-7,-9,-14,-9,-15,11,0,5,0,3,1,-9,
0,7,13,5,3,3,-2,15,7,11,1,-7,-5,2,25,16,10,1,6,8,0,13,11,2,-7,-1,18,4,6,2,13,-2,9,14,-8,3,-5,-2,2,-1,-5,-7,1,2,5,7,6,-7,-9,-3,-4,-2,5,2,-1,-5,-2,10,24,6,-5,-7,-4,0,23,18,11,1,-19,-3,4,2,2,-4,-3,12,-2,-7,-5,3,5,16,17,11,4,-9,-3,3,3,3,2,2,-7,-7,-1,-3,-5,-2,8,-1,6,10,1,-6,4,10,10,14,5,-5,0,4,13,9,-2,-2,8,6,2,10,-3,2,-6,0,12,4,-1,-8,7,-2,-1,9,3,1,1,1,-6,3,-5,-15,-1,12,5,10,0,4,-13,-7,13,11,0,6,3,-3,2,3,11,13,9,9,-13,5,12,9,14,21,3,-16,8,-5,-7,-6,0,5,-9,10,3,-5,6,8,16,10,9,-7,3,4,6,5,-3,1,-7,3,-1,-10,-4,-6,-5,-1,5,-4,3,-2,3,7,-1,9,10,10,4,4,4,22,23,18,-11,-12,-4,10,21,31,2,-1,-10,-12,-14,-13,-22,-12,-3,6,2,-3,-20,-16,-8,-4,11,6,-5,-2,-7,-8,-3,2,-5,-2,2,-4,0,4,-5,1,8,7,5,8,3,-7,-7,13,7,-3,-7,3,19,10,17,2,3,-2,7,19,-3,6,10,3,6,9,6,-4,10,1,-7,-1,-9,-1,-11,4,-1,6,7,4,-9,-7,7,2,2,6,2,-3,4,6,-3,-3,-11,6,6,13,4,5,-23,-22,-3,1,6,-4,-27,-30,-23,-3,-1,-2,-3,-3,6,-1,-6,0,0,3,8,10,0,2,6,-4,-6,8,0,1,5,10,2,-6,0,5,8,4,2,-3,9,12,14,13,-3,-10,-17,18,16,17,6,0,-1,-15,4,6,-3,-13,-3,17,1,-3,-6,-6,8,17,15,6,0,-11,-5,-3,0,1,-8,11,1,-5,0,-2,-8,-9,
3,2,-5,-3,-6,3,-1,-1,-1,3,-1,-6,-6,2,-6,1,-1,3,-6,-6,5,-5,-4,5,2,-2,4,-4,-4,-2,-6,-6,-3,3,-3,6,-1,-7,3,-3,-5,0,6,0,-3,-4,3,1,2,-3,1,-5,5,-1,4,3,-3,2,-5,-2,2,0,-4,-4,-7,-4,2,-5,-5,-3,-1,-4,4,-2,2,-1,2,1,-2,3,-1,-4,-2,4,3,2,-5,-4,-7,5,-6,-1,-4,-4,2,1,-3,2,2,4,5,2,-3,-4,-3,1,-1,-3,1,5,-6,-6,1,-7,4,3,0,5,-4,1,-7,-4,-7,-6,-2,-6,-3,-5,-7,-6,-6,1,-6,-2,-3,0,2,0,2,-6,5,-2,5,-3,-1,-4,-7,2,4,2,1,-2,-5,0,4,3,3,3,5,5,-4,-4,5,-5,-3,-7,2,1,-5,-7,-7,-4,-5,-1,-6,-4,-4,-1,-6,4,-5,-3,-7,1,-5,0,-3,-5,-5,5,-4,3,-7,-2,-3,6,4,-2,5,5,3,-5,-1,0,1,1,3,2,5,1,4,-5,-3,3,0,-3,4,-6,-3,-1,-3,2,-1,-6,3,-1,3,3,-1,3,2,-4,2,5,-4,-3,6,3,-7,-4,-2,-6,-1,4,3,-1,4,1,4,0,2,-5,5,-5,5,-5,5,-7,3,-3,1,-7,1,2,4,-5,5,4,4,-7,4,-1,-4,-4,-4,-6,6,4,-3,4,-2,-2,0,-3,-6,2,1,5,-4,5,3,1,3,4,2,1,5,1,-7,4,4,3,-2,-5,-4,3,3,1,2,2,1,-2,3,-2,1,-1,4,-4,-1,4,-1,6,5,-6,-7,-1,2,-1,-3,2,3,-1,0,5,3,-5,-1,-5,-4,-6,2,-3,6,-3,5,-3,-5,0,6,2,5,5,-4,-3,5,-4,5,4,0,5,1,-6,-5,6,4,1,2,-1,2,4,0,2,3,3,-6,-6,0,1,6,1,5,2,-2,-3,-4,2,6,-2,-6,4,5,-3,
-3,-1,-16,-5,-11,-8,-5,4,14,13,3,2,-4,-8,-5,4,8,-7,-6,1,9,2,3,2,9,3,-2,-5,-1,-2,-4,-2,0,-7,-3,-10,-6,-5,-7,-3,-7,7,7,12,10,5,4,3,16,4,2,5,2,-3,6,4,2,-10,1,-7,-1,0,-6,3,-4,-4,3,-6,0,5,0,-7,-2,4,8,17,10,3,7,17,18,4,-15,-11,-12,-4,-6,-6,-6,-3,-6,7,5,0,-3,-2,6,-1,-2,-12,-1,-7,-14,-6,-11,1,-2,1,4,0,6,3,-3,-4,-3,-3,-9,-3,7,-13,-1,23,18,15,-3,-2,-16,-6,-4,-7,-5,-18,-1,6,7,7,-6,-7,1,9,5,4,14,13,2,0,5,-8,-15,-10,-3,-3,-1,0,3,-8,-9,-4,-10,-14,0,2,-7,7,-6,6,2,2,3,9,16,-3,2,11,28,-5,-7,11,25,7,0,-22,-12,-8,-8,-6,-8,-12,0,3,-2,-5,-8,-3,-1,8,-7,3,5,-5,-5,0,-3,3,8,2,13,10,9,0,-6,-7,-15,-10,-6,7,8,-14,-30,-7,8,-7,1,0,-2,15,14,-1,1,-8,7,9,37,34,0,-15,-16,3,5,3,-6,-14,6,-6,-3,2,-5,-7,-19,-11,-15,-15,-4,7,8,-5,1,-5,12,-2,20,15,-5,-1,0,6,-3,4,9,4,9,-2,2,-6,-14,-20,-15,-2,-14,-2,-19,-4,1,1,-8,16,11,4,11,8,5,2,11,5,0,-1,-12,-7,5,-2,-12,-1,-6,4,-6,4,1,-13,3,-5,9,-10,-5,-3,6,0,27,22,-4,-7,4,5,5,8,-22,-7,3,-11,9,2,0,-24,2,1,-7,4,-2,-1,1,15,13,-7,8,3,-11,-3,-3,3,0,-4,-1,4,7,0,-2,-7,5,-5,-5,-6,-12,-6,7,20,-3,2,20,21,8,-4,0,-10,2,19,20,6,-13,-21,-8,-6,-1,-14,-12,-5,-3,9,13,0,-1,0,8,13,
7,10,16,-6,0,9,2,4,-8,-3,6,6,1,9,-6,0,-4,-4,-9,6,6,-3,0,10,-3,-15,1,12,-14,5,7,15,-10,5,7,-6,-5,4,11,10,9,-2,-17,-8,1,5,-2,-3,0,10,9,0,0,-1,-1,0,3,1,-3,-17,-1,4,8,9,2,-13,-3,8,0,0,-4,-5,-9,-7,-2,3,6,7,-6,-17,-3,7,10,10,0,1,1,1,4,11,2,6,2,11,14,4,-1,-1,7,0,1,5,5,9,8,2,-3,-6,-4,-8,5,6,-3,-3,-5,3,-8,3,-4,9,10,-3,2,-6,-2,9,-2,-9,-3,9,2,10,7,4,-3,13,19,4,11,-1,-4,-19,-17,-13,-2,-4,10,7,15,9,5,21,5,1,3,-10,0,-8,10,11,4,-7,-5,-2,-11,4,-4,5,-10,3,5,1,-1,2,-6,-2,9,-3,3,2,13,14,6,2,17,4,5,7,1,8,8,16,13,7,8,5,9,3,-4,9,10,9,1,-2,1,-10,-8,-3,5,-1,-3,0,-3,-10,-4,2,-1,10,11,0,1,6,3,2,6,-15,-39,-12,15,8,3,-3,-23,-29,4,5,16,2,8,3,10,14,4,-4,1,6,2,6,10,16,16,8,8,-6,-9,-9,-6,-7,-5,1,2,2,2,-14,0,15,-1,4,7,2,-2,1,13,-3,9,27,10,4,2,6,-4,4,7,-3,9,-3,3,5,-9,-9,-11,-12,-1,6,5,0,13,13,3,-4,6,-2,10,15,19,6,11,5,9,-2,13,20,3,1,-10,4,-3,-8,28,-1,-8,-15,-1,-3,0,18,5,5,-8,7,12,21,0,1,-3,0,2,2,-26,-19,-13,-3,4,5,10,7,0,6,8,-2,-13,-9,-3,-6,-1,1,11,-10,-7,-7,-4,-8,4,-1,-5,9,-4,-4,-8,11,13,-2,-1,-5,3,-1,4,15,-1,2,18,18,14,9,5,-20,-5,2,4,7,8,5,
-2,2,6,5,-13,-8,3,10,-3,5,9,4,4,-5,12,10,-1,7,20,6,2,-6,-10,-19,-5,18,-1,-7,-9,-9,-8,16,3,-13,-7,9,7,1,-1,-5,4,-6,6,10,8,4,1,0,-3,-3,-2,-4,2,15,3,1,2,8,15,1,-12,-20,-4,13,31,39,16,-3,-16,-6,-6,17,1,-6,-7,2,11,-3,0,4,5,0,-4,5,0,-1,4,6,-2,4,5,8,3,0,-8,0,3,-2,13,8,7,3,-3,-2,4,7,14,15,11,1,-8,3,-5,8,-3,-4,10,3,-1,-3,0,-5,-7,1,-4,-7,5,-4,5,5,9,-4,6,6,7,-1,3,-2,0,7,-5,9,14,9,6,3,-2,4,3,15,6,1,9,-1,7,7,2,4,8,6,-17,-3,12,5,30,1,-5,-11,-7,-4,-13,-3,-13,-15,6,-4,-6,-10,0,-17,-4,18,6,5,-6,4,4,5,9,3,9,1,1,1,6,-4,5,-5,0,4,-2,4,-3,0,8,3,11,9,0,2,4,17,20,9,-9,-22,0,14,30,33,-5,-14,-12,3,5,8,14,-20,5,20,13,1,7,2,-1,26,28,9,-2,7,5,0,1,2,8,11,-2,0,9,1,-4,-11,8,-9,7,5,11,1,-11,-5,-9,-26,-3,-1,-1,-14,-7,-6,-17,3,9,-11,-10,1,-3,4,11,5,-1,8,0,7,2,-3,-5,6,1,8,15,1,0,9,6,-4,-8,-1,-1,2,2,-3,-6,-7,-5,-25,10,7,-3,14,-6,-7,-46,-17,14,-8,6,-1,-21,-41,-25,2,-4,-4,-1,-9,-11,-2,-5,-1,-1,1,-5,6,4,-1,4,-14,-1,-8,0,12,2,7,-8,0,8,8,9,2,-2,0,3,5,8,15,-6,-2,-29,-2,4,0,29,-5,-15,-9,-16,-8,-17,-3,-7,-11,-9,-2,-8,-2,-4,-12,-8,2,-1,1,-4,-1,-6,8,4,15,5,6,2,-3,2,-7,
-4,-1,-1,-4,4,0,2,24,10,9,-8,-9,7,19,18,2,5,4,0,5,3,-3,-1,6,-5,-8,-8,1,8,-3,-10,-4,-2,0,0,11,1,6,5,10,2,-7,7,4,0,8,0,-7,-14,6,-3,5,2,2,1,6,3,11,-1,1,-14,-3,-6,1,25,7,-4,-2,16,15,7,8,0,3,11,9,6,3,2,-2,-18,6,8,2,9,4,-6,4,6,12,6,1,-4,9,4,11,5,6,7,-4,-7,0,5,4,2,0,13,14,-6,-12,-1,10,1,6,-5,2,2,-3,8,6,4,-6,-2,-7,0,-5,13,-5,4,5,8,12,3,7,-2,9,10,8,-1,-9,1,3,0,4,4,-13,-7,3,-3,2,12,4,4,1,8,13,27,12,-1,4,-9,-2,3,0,-7,-7,-7,22,-1,0,-11,-7,-6,10,13,6,-5,-9,-9,-3,9,5,7,4,4,9,9,2,2,4,5,5,6,2,2,-5,-2,-5,0,-3,0,10,-2,-6,7,-2,-14,-10,4,6,2,9,2,8,0,6,2,13,27,16,13,27,36,15,16,9,-3,9,41,21,4,-1,1,-4,4,3,9,-4,2,-2,2,10,-7,-6,-1,2,21,-7,-4,10,20,12,5,16,8,-12,-6,13,19,-5,-8,-16,3,4,4,4,1,-10,1,1,-14,-4,13,-6,7,13,12,6,10,16,11,-6,9,5,7,-8,-14,-4,1,-1,-4,6,-14,-1,4,-1,4,-11,2,1,7,-5,11,31,19,1,5,2,4,7,1,21,-6,2,-10,4,-20,-28,35,8,2,-11,5,5,-13,20,14,2,-5,-4,1,-6,-9,3,3,-10,5,0,-11,-12,-14,1,-1,7,-4,7,5,7,4,-3,21,26,16,-12,-14,3,18,1,11,9,3,0,11,20,-1,-5,-6,-12,-12,0,0,1,-6,-8,-11,5,14,21,7,5,8,10,15,10,-2,12,-1,2,10,-3,-11,-4,
1,-1,-9,-3,6,4,5,2,4,2,-2,13,1,0,4,-3,2,2,-1,-3,-5,-1,2,6,1,0,-7,-2,6,-1,0,-5,2,7,3,0,2,-9,1,6,0,10,-5,-6,-8,2,-2,8,-4,-5,-2,1,-10,-7,-2,4,4,-14,-8,-6,2,1,8,0,-2,-5,1,-5,7,-3,-3,-2,-8,0,-12,-6,-3,2,3,7,-10,-1,-2,-9,-5,6,-6,2,-2,5,-1,2,-1,-9,8,6,2,-5,-1,1,-1,1,7,1,5,9,5,-1,3,1,-3,-5,2,1,9,3,-6,-4,-9,4,2,-1,-7,1,5,-4,5,0,-4,7,8,7,-4,1,-2,-1,3,5,7,-1,0,-3,-3,5,5,-8,7,-1,-13,-5,-1,-1,0,3,0,5,2,8,-3,-8,4,9,8,7,-2,7,-12,-1,6,6,4,4,2,-7,1,2,0,5,-2,-5,12,-1,-5,4,0,-3,-2,5,-5,8,1,-6,-3,6,10,-3,-2,-1,8,7,7,2,8,2,0,0,-5,-2,1,-4,6,-1,2,-12,-20,-6,-6,-6,5,0,-5,-1,5,4,12,5,-1,3,4,7,-4,6,7,6,-1,-3,-2,-6,-2,1,1,4,-1,3,1,-2,-7,5,3,11,0,-4,-1,4,0,-1,8,5,-2,-1,5,-2,-3,0,0,-1,4,5,1,-9,-7,-9,4,2,5,-1,3,8,3,10,-3,7,-11,4,9,14,2,1,-10,-12,4,4,-2,6,-1,-5,-2,-1,12,-2,-2,5,4,18,-2,10,4,-7,4,9,30,1,2,3,-1,-1,-1,13,10,7,-1,-4,2,2,3,-1,12,-1,9,-6,-5,-2,-10,9,4,8,-5,6,-1,-16,-1,3,2,-2,-8,-3,-1,1,-4,-5,-2,3,-8,1,-2,1,9,0,9,2,0,5,-8,-2,-4,-5,1,-8,-1,-6,-3,-4,8,-5,4,1,3,5,8,-3,-7,-3,4,1,5,-3,-11,-6,-1,-3,-4,-5,
0,1,7,-3,11,9,3,-14,2,6,4,2,-2,-7,-10,4,1,-2,-9,-4,-3,11,-5,3,-2,-1,-7,5,-13,-9,2,1,-1,-1,-1,-10,-14,3,-3,-6,-1,2,-7,-7,-8,-6,1,3,3,1,-3,2,-1,-7,1,-2,-1,-10,-2,20,28,20,1,-3,-10,-1,18,30,18,-2,5,5,-7,1,-2,-1,0,8,5,-10,-1,-7,-9,0,-2,-1,9,5,6,4,-1,-5,-8,4,4,-1,5,-3,-1,9,3,6,5,-1,2,-3,-5,-8,0,10,-2,-14,-1,0,8,0,3,-1,5,0,-1,-2,-1,0,3,-1,-4,-9,8,3,-6,-5,-5,-8,-8,-2,6,1,5,2,-9,-10,-11,-3,11,3,-3,6,6,-4,1,12,4,3,-6,1,-8,-15,-12,-2,20,-2,4,2,7,1,21,10,6,-3,3,-4,-6,6,1,-3,-5,-1,-5,1,-1,-2,-13,-3,9,5,-5,-6,-3,-1,-4,1,-3,-6,-4,1,2,1,2,-6,-2,-2,6,1,1,-3,11,4,-2,-1,-6,-10,-12,16,39,27,13,-8,-9,3,16,23,4,-2,-2,-3,-13,-11,-1,-4,6,-3,-16,-25,-6,-3,-8,0,-5,-2,-1,-5,8,8,-6,-7,-1,14,-1,-6,7,-1,-1,8,11,1,-3,-8,-12,-4,16,20,3,-11,-9,-2,-2,-3,-2,-6,1,-2,8,-6,0,13,12,-2,1,5,-8,-4,-3,-9,-7,-4,14,2,-7,-4,2,3,5,10,3,-2,8,9,-5,-4,-6,2,1,-20,-17,-13,-1,-21,-2,-1,28,-1,-19,-13,-8,-3,7,15,0,6,-7,2,2,2,-15,-15,6,4,-4,5,4,11,7,8,1,-2,-2,0,-11,-5,1,3,7,6,-3,3,1,8,-2,-2,-15,0,-7,5,9,16,10,-2,2,3,5,7,10,12,-1,1,2,7,2,-3,10,-16,-3,-5,5,2,-1,-5,-10,-6,4,3,7,6,6,-18,-9,-3,-2,-5,2,3,
-4,-7,-1,-1,0,-2,-11,0,1,6,-1,-4,8,11,11,6,4,-4,-3,0,-8,2,-4,6,-5,1,-2,-16,3,6,6,-2,1,4,-8,11,9,-3,-6,0,4,4,-1,-4,2,-8,-5,6,5,-9,-1,-2,-10,-3,-3,1,-5,8,22,4,-5,-12,-8,-6,5,11,1,-20,-5,0,-7,6,11,3,7,4,2,-4,6,7,11,2,6,3,-2,1,0,6,-4,-6,1,-5,-10,3,-3,6,3,-5,-3,-3,-4,0,-3,4,-9,-2,6,13,6,4,2,2,2,-4,4,1,-5,-1,-10,-4,-6,14,15,7,11,-10,3,9,-1,-1,6,7,6,-9,2,7,-2,2,-2,6,5,10,4,2,-2,3,7,2,-8,7,4,-15,-8,4,-3,-6,13,13,12,7,-7,-3,5,2,-1,10,-5,0,-7,4,2,5,-4,-12,9,1,-2,3,8,9,5,5,9,3,-1,2,8,5,3,-2,-3,0,1,-1,0,4,-6,0,-5,0,1,3,4,-8,3,1,-1,1,1,4,0,9,5,-7,-12,-16,-10,9,15,6,25,2,0,10,-2,9,15,20,5,10,2,0,12,10,3,5,13,6,-8,-6,-1,-8,-8,-10,-6,-10,-5,-2,1,11,3,-6,-4,0,0,-2,2,-7,4,-4,-9,-11,-10,-5,-4,-8,3,-4,-2,6,12,3,-1,1,6,-8,-7,5,1,11,-2,-3,2,-2,1,9,2,-6,-1,0,9,7,-12,-7,3,2,-3,-12,2,11,-7,-2,3,0,-5,4,1,1,-7,-3,-36,-3,-8,12,-4,-4,8,-26,-5,-5,-5,0,-8,2,-26,-12,2,1,-9,-2,4,-46,-31,-3,-5,-1,-3,-1,-15,-13,-2,-3,-4,0,-2,-1,8,-1,-6,-9,9,-5,3,9,2,1,-4,9,-3,-6,-9,5,-15,9,-8,2,17,12,-1,-6,-4,12,8,13,23,11,7,0,3,1,-6,-11,13,6,10,17,2,4,-3,0,5,15,
9,-1,-3,0,6,11,6,9,2,-6,2,10,-4,-3,-11,-10,10,1,-4,-12,-11,-5,5,4,1,11,-2,3,4,5,-5,4,12,2,0,-1,-5,-4,7,2,-1,-11,3,-5,-10,-7,3,4,0,2,3,11,6,4,12,13,10,9,-5,-8,9,1,13,1,1,2,7,11,16,8,4,-3,-5,2,-16,-10,-2,12,12,7,9,1,0,3,3,-1,10,2,-1,1,10,4,0,-2,-3,-4,3,3,3,0,5,-5,3,1,4,11,0,-5,-2,3,4,-2,-5,3,-7,0,-3,-10,-2,1,5,2,-8,8,1,13,0,-2,4,5,11,1,-2,5,1,-15,-3,1,-1,-2,10,7,8,8,3,11,6,9,7,9,1,7,6,11,9,4,-5,-3,-6,2,5,0,1,-5,-7,-15,4,4,1,0,-5,-2,-3,-4,-10,8,6,3,11,1,-1,5,-7,-6,-6,8,2,9,7,-3,-5,-6,-10,-2,-1,2,10,8,3,5,1,3,6,10,3,-6,-8,-2,-3,4,4,3,2,-5,13,11,6,2,0,-3,16,5,2,4,6,-12,14,5,-14,4,5,9,16,8,-14,6,13,9,12,9,-1,-11,6,4,10,8,-6,-4,-6,-10,1,-1,6,-1,-7,2,8,1,-8,8,4,3,0,9,-2,-6,7,1,5,-5,10,-1,3,6,-6,-1,15,12,-7,-3,7,-1,-9,0,-12,-9,1,4,13,5,4,9,9,7,-4,2,10,4,-3,0,-1,3,3,17,0,8,1,4,-1,11,20,3,9,-8,11,5,2,17,-19,10,2,9,1,3,25,-5,-5,-3,8,0,-10,13,26,4,12,-5,2,-2,39,34,15,8,7,11,6,4,3,8,14,6,4,4,-3,-13,-2,3,6,-10,-6,-16,-9,-5,-8,-15,10,0,-16,-11,-4,-5,-11,-1,-1,9,9,-1,7,-1,-19,-1,1,1,7,-4,-7,1,-6,-17,-8,-5,-1,1,
10,8,-2,2,-11,-10,-1,3,-5,-13,-14,7,13,-1,-13,-20,-3,-8,6,-2,-8,-10,9,-2,3,2,-14,-14,9,6,-1,18,12,-4,6,6,6,5,2,-6,-8,4,0,2,-3,-7,-9,-5,-8,7,9,14,5,12,11,4,12,7,-3,-6,-17,1,8,13,4,-8,-20,-12,-2,10,5,0,-1,1,-20,-11,8,9,10,0,3,7,19,17,5,3,-1,8,9,11,10,10,1,-4,-3,0,2,11,5,-3,2,-4,0,-4,5,6,-9,-6,-14,-5,1,9,3,-1,-5,-6,-1,-5,-5,11,10,3,9,1,-4,11,2,6,2,15,16,1,12,2,-8,-5,-4,-6,4,4,1,-20,-6,-6,-2,1,8,10,6,5,0,5,3,2,11,10,13,15,-6,-9,-11,-8,-6,-4,-14,-18,-17,7,-1,-2,-6,1,-11,-18,-7,6,11,13,5,-4,7,23,11,5,-4,8,0,10,7,8,4,4,-13,-4,-5,-1,7,11,8,5,10,3,7,4,1,-5,-16,-5,-4,10,1,9,-5,-4,-2,0,8,14,25,17,26,-5,-1,9,2,-2,2,5,6,15,10,4,3,-3,-24,5,14,8,13,11,10,16,2,-1,12,12,-9,0,1,6,-3,5,6,-20,-14,-7,-4,8,-2,-1,-21,-8,2,15,-5,-24,2,-1,9,5,8,-17,2,2,9,9,10,7,-3,7,9,-9,-9,9,-8,3,3,3,-1,-7,-6,3,-12,15,-2,-1,0,4,9,1,3,7,7,29,35,9,1,3,3,5,15,42,26,8,2,-1,-12,-15,26,5,-1,-2,0,0,16,12,0,1,3,4,-2,21,17,2,9,3,7,8,16,13,-4,-2,6,14,10,-2,4,3,2,7,-10,-4,-1,-17,-20,-1,14,-14,-5,-9,-8,-13,-8,-3,-1,-5,1,-4,-19,-15,-3,7,-3,-4,-3,6,3,25,-1,-4,-8,-1,4,10,11,-9,-8,1,3,6,5,3,
1,-9,-4,5,4,4,-2,-14,-1,7,2,1,-3,7,7,8,-5,-11,-6,-1,5,8,-8,-15,3,12,-12,-6,2,-2,-7,15,2,-14,-5,8,10,-4,0,-7,9,13,-2,1,-2,-3,-1,16,15,-6,4,4,-2,-4,-5,0,-1,0,12,12,12,-2,2,3,0,8,0,-3,-8,-4,4,25,23,1,15,20,13,2,2,8,23,6,-6,11,-2,5,-2,1,-9,-7,-1,-6,0,0,0,7,9,0,-4,-8,4,5,1,8,1,-5,4,11,0,-1,3,0,-2,6,-4,2,-10,2,3,4,4,7,25,13,-4,-3,11,15,-7,5,0,-6,4,-2,5,8,-2,-2,16,7,6,7,1,1,3,10,7,-9,-2,3,8,-8,-2,-2,-8,-8,-6,1,10,9,9,1,3,4,5,-4,-10,11,3,0,7,16,-8,-11,25,-1,-4,-1,26,5,-3,18,-2,8,0,-7,-1,12,10,-1,8,3,-11,11,8,3,1,-10,-4,-1,3,6,-5,-2,-1,7,-3,2,-3,1,0,5,9,1,-2,-6,0,8,6,15,24,1,4,7,10,29,11,-15,25,27,19,1,1,0,-11,15,10,8,-5,-7,7,6,1,3,0,-4,-7,1,12,17,6,-3,-2,-4,-1,5,-12,-6,5,-7,-7,1,-3,-5,-6,-6,-5,-8,-16,13,14,-12,-4,9,1,-4,4,-2,-4,11,1,1,0,-6,-7,10,16,-8,2,-4,6,6,5,0,-5,2,-12,-19,-6,1,-1,-6,-6,-15,0,-10,-7,-5,-5,-20,-28,1,-9,-2,-7,0,-3,-6,-11,-10,-16,-5,-2,-23,-20,-16,4,-2,-3,3,-8,-12,-10,1,5,-1,-1,-7,-22,-11,5,3,-7,-8,-2,-5,5,1,-4,-5,-7,-6,7,12,6,12,5,5,-3,6,-2,-7,-1,11,0,-3,15,15,0,-13,9,3,-7,10,26,-1,-7,1,5,13,-6,-6,10,11,12,-4,-3,-1,-2,8,12,15,
6,1,-5,0,-1,-6,6,2,6,-2,-2,3,6,7,1,6,-7,3,7,-1,3,8,3,-3,13,9,2,3,-3,-5,-9,0,-3,-10,-1,2,4,-11,-8,1,-9,2,-3,5,11,8,7,8,-4,5,10,11,8,3,8,5,1,-2,-11,0,-2,6,3,4,2,3,-5,5,3,9,3,12,-2,-1,5,1,5,1,8,13,-3,3,-13,-5,0,4,1,-7,-3,-3,1,8,11,4,0,3,2,4,6,3,10,5,-3,-1,9,4,0,-2,0,10,4,13,1,3,5,10,14,4,11,-1,10,-6,-3,-1,-3,-2,7,-1,0,-1,-8,-9,3,1,8,2,8,-1,3,-1,-4,1,8,17,16,3,-1,4,-5,-10,8,2,1,1,7,6,1,2,-4,-9,7,-1,1,9,12,-3,9,18,0,8,19,18,8,1,10,-2,-7,-6,-1,3,-1,-10,0,2,-3,0,-7,-4,-2,4,5,0,3,6,7,-1,2,1,3,10,-3,-2,11,5,9,12,5,12,6,11,5,-6,-5,18,-4,-2,11,2,-4,0,-26,-14,10,5,8,22,18,-7,8,2,4,6,17,14,3,-10,-24,-9,1,2,-8,-9,6,11,7,7,-9,-1,-1,-9,-10,-8,7,11,7,6,1,14,12,10,11,16,22,7,-1,13,11,-8,-6,-3,-6,-14,-8,-1,-1,-5,-6,-7,-10,-7,1,-2,9,7,6,10,1,7,1,11,17,1,5,4,-2,0,-8,3,1,-6,-6,-4,-6,-14,-3,-10,1,3,3,3,19,1,2,0,-11,3,9,32,12,15,5,5,-7,2,3,3,1,6,13,2,0,10,13,-6,3,-3,-2,0,12,12,5,0,-1,-1,2,0,2,10,1,10,-7,-5,-6,-4,6,-1,1,5,9,7,18,9,9,16,5,6,18,11,4,0,0,-4,0,4,-6,-9,-12,-14,6,6,-6,-3,-11,-16,-10,-13,8,12,8,2,-1,-3,
-4,-1,-10,-3,-1,4,5,-14,-4,-4,-7,-9,-2,0,1,4,2,4,-2,0,1,-2,-4,2,5,-4,10,2,-2,2,9,8,2,-4,4,-4,-6,0,6,-6,-11,4,-11,-14,-13,-4,-8,2,2,-6,2,-3,11,-3,-6,-2,-5,-2,12,17,26,4,7,2,-11,7,8,4,-3,-8,7,0,-9,-11,-7,3,-6,2,8,10,2,-6,0,-2,-2,5,12,12,7,-4,1,4,-2,0,-3,-11,-7,-5,-1,-11,-17,-9,7,10,1,-3,-3,-4,-7,-3,8,5,-2,3,-5,0,-6,-5,-4,2,5,6,3,7,-1,7,-3,1,13,2,-5,-2,-3,-3,-4,-6,1,-6,-2,7,4,10,-3,-4,-4,-2,-3,0,-7,-3,14,-6,7,1,3,-13,-46,-7,9,15,9,6,-7,-3,10,10,12,-4,10,1,-2,-4,4,-8,-5,3,8,7,2,9,3,10,-6,2,4,8,9,-1,3,-1,-5,-1,-9,-12,-7,1,-6,-6,-13,-10,1,0,-2,-5,0,4,8,6,0,8,8,5,10,25,2,-4,-3,3,-9,-2,-5,6,-13,-6,-6,-1,-5,6,3,-17,-1,-6,3,9,-2,1,2,-6,6,2,22,24,11,2,3,0,-11,-18,-11,-2,4,3,-5,1,-13,-7,-11,5,1,-3,5,4,-9,-7,-1,5,11,8,-2,-1,5,10,10,-2,-8,-6,-5,6,-9,1,4,-10,0,-2,-4,-2,2,-2,-5,-1,5,-9,-1,0,-6,-4,-4,-17,-3,4,-2,0,-6,-12,-8,-4,-2,5,2,-15,-14,-6,-11,-2,6,-4,16,8,5,-1,2,-3,6,8,-8,-1,0,1,1,-2,1,-19,-14,1,-7,-3,-5,5,-12,-7,1,-2,6,-3,-3,-1,6,-1,3,-2,0,-15,-22,-11,4,13,1,1,4,9,-1,8,7,-3,8,5,8,-2,4,-2,0,3,5,13,8,-9,3,4,1,-5,10,3,2,1,14,-12,-12,-13,-13,-16,-7,-4,
0,3,-4,-2,-1,-6,0,5,-1,1,1,-3,0,0,0,4,-6,1,0,-2,2,-2,3,-2,-5,-7,-6,-1,5,-4,4,-6,-7,3,-4,-3,-3,1,0,-4,-6,-6,5,2,-7,-4,5,-1,-4,-5,-7,-2,3,4,-6,-3,0,-4,1,-6,-1,6,1,-5,-4,-6,5,-6,6,-3,1,3,3,-2,3,-6,-5,-2,1,0,-3,-1,-6,-3,5,-4,-4,2,-7,1,2,-6,-7,3,5,3,-3,-2,6,0,3,0,-1,0,0,3,6,5,-6,-2,-3,3,0,1,3,-6,-3,-6,-4,-5,1,2,-1,2,5,6,-3,2,-5,-1,3,-7,-3,-5,-5,1,-2,6,4,4,-6,3,-2,-6,4,-5,-2,-5,3,0,6,-1,3,2,1,-2,1,-5,5,2,2,1,-2,5,-6,1,4,4,-7,-3,2,-7,4,-4,0,2,5,-3,1,3,6,6,3,1,-4,3,0,3,6,-2,0,-6,-6,4,-5,6,6,-3,-5,-2,2,-7,2,2,-5,-1,-5,1,0,5,3,5,-5,-3,-4,0,1,0,4,-4,-5,-6,0,-5,-1,6,1,3,-7,3,-4,-2,4,-5,-4,4,4,6,-2,-3,-4,6,4,4,4,5,2,-2,3,0,5,2,-4,-5,-1,5,2,-7,6,-2,5,3,0,-1,0,2,-2,-5,4,0,-4,1,3,-6,-2,-2,5,-5,-3,5,-6,5,3,4,0,2,-2,2,-1,-5,3,-6,-6,-2,2,-1,4,-6,4,-7,-5,-6,6,5,3,5,4,3,-5,2,2,3,-3,1,-6,1,4,5,0,-5,0,4,3,-4,-3,1,5,-1,0,4,-1,-6,5,-4,-3,0,-5,5,6,-1,-2,0,0,-5,-6,2,2,3,3,1,-1,-4,-3,3,-1,0,-1,-5,-3,-5,2,-1,5,-1,-1,-2,5,0,-2,-6,5,4,-5,-2,-5,3,3,-6,-3,0,-6,-1,-5,-5,3,-2,-2,-6,-2,0,-3,1,
5,3,3,-5,1,0,3,-11,-3,0,3,1,-2,-2,-14,-10,8,3,-6,-8,0,-12,6,11,-7,-6,8,-2,-5,9,-2,-9,7,9,1,-4,2,10,-6,-2,1,6,-6,1,0,5,4,0,11,0,6,2,6,2,5,5,1,-13,-14,14,17,16,14,-2,-21,-24,1,13,14,6,3,-16,-10,0,-2,-14,2,3,4,1,-1,-12,-13,3,2,1,6,5,0,-5,-5,-3,2,-1,0,-3,5,6,-2,-1,5,-1,-4,-3,1,-2,-5,-1,-2,8,8,4,-2,-15,7,8,-4,1,-2,-5,-4,8,4,2,11,-3,5,10,9,-7,-7,-2,6,-2,-7,4,2,-2,2,6,7,-5,0,-3,5,9,10,2,-3,-10,-2,-4,3,0,-1,3,2,-9,-4,-5,20,-7,-7,4,-9,4,13,10,-2,11,10,5,6,4,-7,5,13,4,-2,-4,-5,-18,-9,1,-2,-3,0,-9,1,-1,-7,3,4,-9,-1,7,4,10,12,-1,1,-8,9,-2,-10,5,8,13,1,5,-1,-22,-21,-7,19,22,9,-9,-35,-29,7,0,2,6,6,-2,9,23,-16,-25,-4,1,5,10,0,-10,-10,9,7,3,-10,-3,11,2,5,1,-8,6,-9,-8,-16,8,-2,-2,9,1,5,-3,3,3,19,12,0,-4,-7,1,2,11,5,-12,-8,-2,6,-9,-1,-14,-11,5,-6,0,-7,3,-5,5,-4,4,19,0,-4,10,4,7,7,10,-3,0,-1,-3,4,-5,-2,1,-1,5,-11,1,1,-6,-2,2,37,7,-4,11,3,1,15,32,13,4,16,8,9,-1,7,1,-2,1,2,4,-8,-4,0,2,1,12,1,5,16,26,10,5,8,4,-4,-9,-4,-2,-2,1,-6,2,-3,2,10,10,7,-6,-7,-5,5,6,15,14,4,10,6,5,9,-3,-7,3,17,5,3,0,-5,-4,-6,2,0,1,-9,-9,0,0,-2,-9,-5,-3,-4,12,
4,1,-2,3,3,-4,-7,-4,6,5,-4,-1,1,-1,-1,-3,4,4,-4,-4,-5,-5,0,3,4,6,-1,-4,-7,-5,-7,-2,0,1,1,1,0,-1,-1,4,1,2,2,6,4,0,-5,-2,2,4,-5,5,-6,-2,1,1,-2,-4,-5,-2,-3,-3,4,-1,0,-3,5,-6,-1,-5,1,4,3,-7,-2,-5,1,0,6,-5,1,4,-6,-3,-3,5,5,-2,4,1,-5,-6,-1,4,-6,3,0,-3,-2,-2,4,4,2,-6,5,-7,3,-6,-3,5,0,-4,-4,-1,-6,5,-6,-6,0,0,-4,-4,5,-6,2,1,2,-5,1,5,3,-4,0,6,-1,4,-5,-4,4,-7,-5,2,4,3,3,-3,-7,0,-2,0,2,-3,0,-3,-1,-6,-3,1,1,6,-4,-3,-6,-7,3,-5,5,-5,-3,5,-3,2,-3,-5,-7,5,1,2,-2,6,-4,6,-4,2,-6,-4,-2,-2,-2,-7,6,2,1,1,0,2,1,-4,2,-3,3,3,-4,0,-7,3,-2,-6,0,6,2,-5,3,-6,5,-5,4,5,-5,0,-4,2,-6,5,1,-4,-1,3,-7,-3,0,-6,0,-4,3,2,-7,-3,0,-7,-4,-3,-1,1,-5,2,-2,6,-2,1,1,-1,-6,2,0,4,-3,3,5,0,-3,0,0,1,5,-6,-2,5,-3,-5,3,5,0,0,3,-1,-2,-6,-2,4,4,-4,-2,-2,-5,1,-4,-6,-1,-5,-4,-2,3,3,-5,-5,6,6,2,0,-5,1,0,-3,-3,5,2,-2,-2,4,-3,-1,4,-6,-2,6,-4,-7,-3,-4,-3,0,1,1,3,7,-6,-2,6,3,3,0,-1,3,6,1,-3,-4,-5,1,3,-5,-5,5,2,-3,-6,3,-5,4,2,-4,-5,-3,3,3,3,2,2,1,-7,4,-1,-4,-1,0,-6,-2,-3,-4,-4,0,0,-6,-5,0,5,-1,-4,-1,6,1,-7,-3,3,4,5,2,0,4,0,-3,
3,3,-1,2,13,9,4,-3,7,6,-3,5,5,-13,0,11,-9,-1,-2,3,4,6,-3,-6,18,7,-13,2,13,2,-2,1,-7,-2,3,8,-4,-5,-3,-3,-2,6,-7,-9,1,-1,0,5,7,-2,-4,-6,-3,-5,-6,3,6,-9,-5,-7,7,13,8,3,4,1,-9,-4,18,-6,0,6,-2,4,21,5,-2,9,2,-4,4,-10,-16,-9,3,5,5,6,3,-4,-9,-7,-6,0,11,9,3,-5,3,4,6,6,9,5,4,4,-1,-3,8,3,-5,-6,5,3,-2,2,5,5,1,0,5,-1,13,6,-7,-6,6,16,-3,3,-3,2,4,-12,9,7,7,-1,-5,0,6,15,25,13,4,-1,5,-2,-8,3,7,9,-6,-3,1,5,-3,1,-14,2,14,0,-5,7,3,-9,0,3,11,-1,3,10,2,11,6,5,6,-4,8,4,-5,-17,-3,2,-2,-2,4,-7,-2,-7,-9,-5,-5,-4,4,0,-2,2,-1,-3,1,2,4,-4,0,1,-5,-8,-3,-7,-2,-14,-3,-2,9,14,2,-3,-8,-17,-20,15,18,1,0,13,6,-5,4,0,-7,-3,12,15,13,-15,-25,-6,1,2,20,13,-4,-6,-2,-3,6,6,9,9,0,2,4,9,-3,6,-1,5,-5,-1,9,-5,2,7,-2,4,9,-7,-6,6,-1,-8,2,7,-6,-11,2,-17,7,6,0,-6,-9,-8,12,2,-3,-4,3,-1,16,2,13,7,-5,4,1,3,4,-1,-5,5,-12,-11,-14,-9,-13,-14,3,-9,-7,-27,-14,-5,1,-8,20,26,-32,8,-8,9,-4,5,-4,-10,15,7,-2,5,-4,-25,-17,-4,-3,2,-1,-5,-28,-16,-6,1,-1,1,-8,2,1,-5,-3,-5,-5,-5,-8,-2,2,2,3,0,-4,2,-1,1,7,11,14,1,5,20,19,6,-8,8,1,11,10,1,-13,-9,4,13,5,5,0,-7,-5,7,-1,1,-3,-8,-4,3,
4,0,-2,-8,7,6,7,3,1,-5,2,-2,-4,2,-13,-7,7,1,-1,-10,5,-2,2,12,-1,-1,4,5,3,-1,1,-4,12,15,6,-15,-1,2,2,4,-2,-8,-6,-11,4,0,-3,0,6,-1,-5,6,7,2,-1,8,7,-10,2,-4,11,12,10,-3,-3,-17,-3,2,16,5,2,-6,-9,3,-1,-8,-1,-2,12,7,5,-5,-4,-1,-1,3,4,1,1,4,2,-6,-5,-5,-4,-1,-4,6,-3,-1,2,3,5,6,-4,-5,4,-5,-3,-4,6,-7,-2,0,4,-1,2,4,7,2,-1,7,3,13,14,2,-2,7,6,0,5,8,-2,-2,-6,-12,-1,-3,-7,-6,11,7,1,8,6,12,5,8,0,7,2,5,-7,4,4,11,-2,-11,-6,-8,8,-3,0,-10,-12,-3,-1,16,1,3,-2,-2,1,3,0,0,15,2,3,1,-5,1,-2,0,-2,-3,1,4,-5,-1,-13,-8,-4,1,-4,5,-3,1,-5,0,-3,2,0,-4,-1,2,-1,-1,-5,5,-7,-12,-7,-4,16,14,17,-4,-3,-21,17,14,6,9,1,-1,15,22,-21,-10,-2,0,18,10,-5,-10,-5,3,-3,2,-1,-10,5,0,3,5,-2,-5,-9,-5,6,10,3,2,4,5,-8,0,-7,-1,4,10,-3,12,4,-2,-3,2,11,2,5,3,0,-2,0,-5,3,10,1,-9,1,-8,-7,5,-4,-5,-6,-1,6,7,3,0,6,13,7,-6,3,-1,-5,2,4,7,2,10,-2,7,-1,-2,-1,14,11,1,-11,0,9,1,14,14,-17,4,0,13,4,-5,10,-9,-5,-8,1,-1,-1,-15,2,4,-2,8,0,-3,14,17,21,6,-3,5,-5,0,1,1,2,-4,4,6,1,-3,-4,3,8,-5,-8,-2,-9,0,3,-2,11,-1,2,0,9,9,-4,-4,7,9,8,10,6,0,-21,0,3,0,-4,-3,-8,3,-10,-3,-2,-3,0,-2,
-3,4,7,-3,5,4,6,0,-2,11,8,3,7,14,-15,1,-6,-2,-8,-5,12,-2,-5,0,10,2,-9,3,0,-7,2,2,2,-2,-8,-5,-4,1,-1,-3,3,3,-18,-1,1,4,4,-6,2,-1,-6,-4,-2,-4,-5,0,-5,-3,-13,-14,-3,22,12,-1,-8,-16,-7,2,30,12,2,-7,-3,-4,10,5,8,-3,7,-9,1,11,-9,-8,-5,0,-7,1,-7,-10,1,2,-7,-3,8,7,4,5,2,6,1,5,-3,5,4,-4,5,4,-9,-3,5,13,-3,-1,6,5,-7,5,6,5,0,5,11,5,3,-7,-3,1,-4,4,-3,0,-3,-4,-7,7,12,11,-3,0,-15,-18,-1,0,-8,-8,12,-6,-9,-2,0,7,4,-2,-2,3,1,-10,-4,7,17,3,0,6,-15,-5,0,24,0,-4,13,10,3,13,-4,-2,1,4,8,14,8,-10,-3,3,2,0,5,-7,-10,-14,0,2,7,3,7,-1,5,9,6,6,-3,-7,-3,-3,4,-2,-6,-7,5,1,-8,-24,-25,-5,3,15,4,-1,-16,-17,0,17,11,-7,4,2,-6,-6,6,10,-1,-1,-9,-20,-13,-18,-24,2,2,-3,6,-16,4,-1,2,3,9,8,-3,0,6,10,4,12,6,-3,-13,-6,17,-4,4,9,5,-4,-2,-2,-6,-5,-2,2,0,-8,-4,0,-3,1,8,-9,-6,-10,-5,1,-3,-3,3,6,-1,-6,-5,-2,-5,-7,-7,-1,7,4,3,10,5,-9,-2,3,3,18,-6,-2,-2,-13,4,-1,32,17,-15,-8,-12,-2,12,30,7,0,-2,-1,4,-6,8,1,16,4,3,-2,-9,10,13,-2,-10,6,6,-2,-21,-18,-3,-9,9,0,-7,-1,-8,5,6,3,1,1,-7,-10,-6,9,28,-5,-1,6,-18,-7,14,14,-2,5,14,16,10,2,-8,-7,2,-7,13,1,-3,-10,-10,-3,4,8,-1,-9,-3,-22,-8,11,11,4,-2,-4,
4,-2,6,1,8,-10,-1,-3,-2,-9,-15,-17,-12,-6,2,2,-5,6,7,7,9,2,10,11,4,-2,-5,8,15,11,-3,1,-4,-2,-2,2,-3,-7,-8,5,2,0,0,-8,-2,1,0,-7,-7,2,-1,3,-1,4,2,4,-1,-3,4,10,15,6,6,3,-1,-16,-5,12,7,10,4,7,5,6,6,10,9,8,18,8,-2,-2,5,4,5,4,4,7,4,-5,-1,-1,-9,3,-5,-6,2,5,4,-2,-7,5,-8,-10,2,3,-6,-15,-18,-12,-8,-1,1,5,5,7,11,13,9,15,3,-7,0,-5,-1,4,12,5,-5,-3,0,8,6,-2,-8,3,-9,-3,-4,0,-3,1,4,1,4,0,3,-1,14,7,1,-2,-2,7,-2,6,0,-5,-10,-18,-3,1,4,-6,-13,3,4,9,4,2,3,4,7,8,20,7,11,-1,-8,-1,-3,12,-4,4,-11,-4,0,0,-1,-6,-4,-5,-2,2,-8,0,5,-6,-1,-6,-3,-10,-6,1,1,-9,-8,-9,-5,3,2,8,17,20,31,24,23,11,16,2,-3,18,24,8,8,19,-3,-3,2,9,-4,3,10,20,18,10,2,-1,4,-1,7,16,-3,-5,1,6,-5,1,-1,-4,-14,-6,-2,3,-7,-8,-9,-10,-8,6,-2,-9,9,2,10,12,9,4,13,4,-1,-6,8,-2,2,6,-4,-1,2,-2,4,-2,-5,-3,6,-6,-9,2,-4,-11,1,7,-1,3,0,-8,4,0,-2,-6,-2,-5,5,14,-7,-3,-2,-11,-1,7,7,13,-15,0,3,-1,-9,-20,20,6,7,-6,-3,-6,-6,1,-4,-1,0,6,3,2,-11,-1,4,-2,-7,5,1,-15,-8,1,0,5,0,-1,11,-2,0,1,4,2,-12,-14,-16,-18,-10,-3,-2,-1,-2,10,5,14,0,6,6,9,-6,4,11,11,0,0,-3,1,2,9,-13,4,-7,2,-10,-13,-13,-2,-1,1,10,6,-2,0,
-5,-1,-1,1,-1,2,7,-8,-3,-3,10,-1,5,2,-9,-6,0,0,-6,2,5,-10,0,18,-7,-22,5,10,-5,7,11,-7,-1,3,15,-3,6,9,-4,4,6,15,-13,-6,3,2,2,0,23,3,-7,-6,1,-3,5,-3,-8,-11,-7,5,8,13,1,-6,-31,-19,10,13,1,5,-6,-10,-15,2,-5,-11,-7,3,-2,1,-7,-11,0,-1,-7,10,7,3,9,-3,-8,-1,0,6,-4,6,3,-4,-9,4,7,-3,-7,2,-3,-2,-18,-8,10,12,2,1,1,-18,-2,-1,-18,0,-1,-9,8,20,4,-11,2,6,-2,0,10,5,3,4,5,0,-7,12,6,5,0,12,1,-9,-15,-14,-13,-1,13,4,8,0,-1,-2,2,-3,-8,-7,-8,5,3,7,9,6,-17,7,-3,21,12,13,-5,0,13,-14,1,3,11,-2,13,10,-1,9,-2,4,-5,11,10,0,0,-2,5,-9,-1,2,6,-1,5,5,-8,6,3,3,-7,-10,-1,3,-11,-2,3,8,0,2,-9,-20,-16,-16,13,18,0,-10,-13,-14,20,10,-12,-2,7,-12,-9,15,-2,-17,-11,-12,-22,6,19,-7,-3,-4,-3,-3,-8,1,7,4,-4,0,-7,4,-3,3,-7,-3,-2,2,0,1,1,7,2,-12,10,12,1,-18,-3,17,-10,20,17,-7,-12,8,13,-2,9,10,-15,9,5,18,0,8,5,-5,11,-4,16,-3,-18,-7,-1,-10,5,9,4,4,-4,0,3,-2,-3,-1,-1,-6,-16,-4,-3,-17,2,2,22,10,-2,5,-15,2,16,1,32,-5,8,-3,2,1,-14,2,2,-6,0,6,12,-15,-17,-5,-6,5,3,3,-20,-10,5,-3,3,0,-5,-8,-9,2,-3,-2,-8,-9,-1,2,8,1,14,-9,-13,-3,0,13,7,18,5,7,10,-5,5,10,13,2,24,11,-3,2,16,15,6,4,11,7,6,3,19,-15,-10,0,-1,-1,4,16,
-5,6,0,7,2,7,-4,-5,10,0,10,5,-9,-10,-7,4,-7,12,4,-6,-9,1,-8,-4,6,3,-14,2,-1,-13,-5,-7,-4,3,3,4,3,2,3,9,13,9,-2,-3,-5,6,11,15,16,-6,-5,-2,6,-3,-5,-5,-7,-10,4,-2,21,10,-2,-10,-2,2,4,22,8,-4,0,-7,-6,9,8,-7,2,-4,4,5,10,-19,-20,-9,1,15,15,2,6,-5,-4,2,-2,3,9,3,5,3,6,-3,4,1,5,8,-2,4,2,1,12,2,3,-2,7,-8,-3,1,-3,-14,-2,-1,-10,3,10,8,-6,-8,-1,10,-5,-6,-9,6,0,-2,7,10,3,4,11,6,14,8,-2,-4,5,0,1,2,6,2,8,0,-1,-2,-6,-6,-11,1,-6,-12,4,1,-8,1,3,-13,12,5,5,1,1,6,1,-2,6,-3,1,9,2,-3,-13,-16,-4,8,-2,-4,-5,-1,-2,0,-2,2,4,4,0,1,-8,0,2,-3,-1,-5,-3,4,4,3,2,-1,1,-3,-2,-9,-3,4,20,9,5,-11,-16,-14,-1,26,13,9,2,12,25,22,2,-16,-9,4,34,45,29,2,-19,-8,3,1,16,17,7,-3,-8,-1,6,8,5,6,7,-6,-5,4,-4,-1,-1,0,3,2,5,-7,8,0,-12,1,6,-6,0,0,-9,-8,6,-7,-3,-13,-13,-10,17,9,0,-4,-4,10,8,1,9,-7,-2,9,0,10,9,14,1,-5,3,-15,-15,-2,-2,-1,-7,-26,-9,-7,-6,-2,3,-13,-19,-27,-5,-12,2,1,22,7,-4,-4,4,4,3,14,-18,-8,3,-5,0,5,-3,-47,-22,-13,-8,8,0,3,-13,-9,-2,0,-4,-1,3,-3,3,0,4,-1,-7,-3,4,5,1,13,-4,4,-11,-3,4,10,4,13,-12,-11,13,20,21,-8,-13,6,-5,8,3,-12,-14,-9,1,7,13,9,5,5,9,7,-4,-5,3,-4,2,8
    );

    constant FC1_B_INT: integer_vector(0 to FC1_N-1) := (
2,-2,-2,0,0,-11,-2,-2,11,4,5,-2,10,0,-2,-4,7,-4,6,10,-4,2,0,2,1,5,1,3,1,1,-2,1
    );

constant FC1_W: mem_t(0 to FC1_M-1)(FC1_N*FC1_DTW-1 downto 0);
constant FC1_B: mem_t(0 to FC1_N/FC1_P-1)(FC1_P*FC1_DTW-1 downto 0);

end package;

package body fc1_rom is
    -- with change ColRow
    function intv_to_mem(intv: integer_vector; constant DTW,P,M: positive) return mem_t is
        variable slv: std_logic_vector(P*DTW-1 downto 0);
        variable ret: mem_t(0 to intv'length/P-1)(P*DTW-1 downto 0);
    begin
        for i in ret'range loop
            for pp in 0 to P-1 loop
                slv((pp+1)*DTW-1 downto pp*DTW) := std_logic_vector(to_signed(intv(M*pp+i), DTW));
            end loop;
            ret(i) := slv;
        end loop;
        return ret;
    end function;

    constant FC1_W: mem_t(0 to FC1_M-1)(FC1_N*FC1_DTW-1 downto 0) := intv_to_mem(FC1_W_INT, FC1_DTW, FC1_N, FC1_M);
    -- constant FC1_B: mem_t(0 to FC1_N/FC1_P-1)(FC1_P*FC1_DTW-1 downto 0) := (others=>(others=>'0'));
    constant FC1_B: mem_t(0 to FC1_N/FC1_P-1)(FC1_P*FC1_DTW-1 downto 0) := intv_to_mem(FC1_B_INT, FC1_DTW, FC1_P, 1);

end package body;
